magic
tech sky130A
timestamp 1624082099
<< psubdiff >>
rect -10 4905 275 4925
rect 515 4905 11800 4925
rect -10 4865 10 4905
rect 11780 4865 11800 4905
<< locali >>
rect 380 6220 395 6470
rect 415 6220 430 6470
rect 290 5820 305 6080
rect 325 5820 340 6080
rect -10 4905 275 4925
rect 515 4905 11800 4925
rect -10 4865 10 4905
rect 11780 4865 11800 4905
rect 1270 4375 1295 4395
rect 1315 4375 1340 4395
rect 1810 4375 1835 4395
rect 1855 4375 1880 4395
rect 1990 4375 2015 4395
rect 2035 4375 2060 4395
rect 2530 4375 2555 4395
rect 2575 4375 2600 4395
rect 2620 4375 2690 4395
rect 2710 4375 2735 4395
rect 2755 4375 2780 4395
rect 3250 4375 3275 4395
rect 3295 4375 3320 4395
rect 3340 4375 3410 4395
rect 3430 4375 3455 4395
rect 3475 4375 3500 4395
rect 3970 4375 3995 4395
rect 4015 4375 4040 4395
rect 4060 4375 4130 4395
rect 4150 4375 4175 4395
rect 4195 4375 4220 4395
rect 7570 4375 7595 4395
rect 7615 4375 7640 4395
rect 7660 4375 7730 4395
rect 7750 4375 7775 4395
rect 7795 4375 7820 4395
rect 8290 4375 8315 4395
rect 8335 4375 8360 4395
rect 8380 4375 8450 4395
rect 8470 4375 8495 4395
rect 8515 4375 8540 4395
rect 9010 4375 9035 4395
rect 9055 4375 9080 4395
rect 9100 4375 9170 4395
rect 9190 4375 9215 4395
rect 9235 4375 9260 4395
rect 9730 4375 9755 4395
rect 9775 4375 9800 4395
rect 9820 4375 9890 4395
rect 9910 4375 9935 4395
rect 9955 4375 9980 4395
rect 10450 4375 10475 4395
rect 10495 4375 10520 4395
rect 10540 4375 10610 4395
rect 10630 4375 10655 4395
rect 10675 4375 10700 4395
<< viali >>
rect 395 6220 415 6470
rect 305 5820 325 6080
rect 1295 4375 1315 4395
rect 1835 4375 1855 4395
rect 2015 4375 2035 4395
rect 2510 4375 2530 4395
rect 2555 4375 2575 4395
rect 2600 4375 2620 4395
rect 2690 4375 2710 4395
rect 2735 4375 2755 4395
rect 2780 4375 2800 4395
rect 3230 4375 3250 4395
rect 3275 4375 3295 4395
rect 3320 4375 3340 4395
rect 3410 4375 3430 4395
rect 3455 4375 3475 4395
rect 3500 4375 3520 4395
rect 3950 4375 3970 4395
rect 3995 4375 4015 4395
rect 4040 4375 4060 4395
rect 4130 4375 4150 4395
rect 4175 4375 4195 4395
rect 4220 4375 4240 4395
rect 7550 4375 7570 4395
rect 7595 4375 7615 4395
rect 7640 4375 7660 4395
rect 7730 4375 7750 4395
rect 7775 4375 7795 4395
rect 7820 4375 7840 4395
rect 8270 4375 8290 4395
rect 8315 4375 8335 4395
rect 8360 4375 8380 4395
rect 8450 4375 8470 4395
rect 8495 4375 8515 4395
rect 8540 4375 8560 4395
rect 8990 4375 9010 4395
rect 9035 4375 9055 4395
rect 9080 4375 9100 4395
rect 9170 4375 9190 4395
rect 9215 4375 9235 4395
rect 9260 4375 9280 4395
rect 9710 4375 9730 4395
rect 9755 4375 9775 4395
rect 9800 4375 9820 4395
rect 9890 4375 9910 4395
rect 9935 4375 9955 4395
rect 9980 4375 10000 4395
rect 10430 4375 10450 4395
rect 10475 4375 10495 4395
rect 10520 4375 10540 4395
rect 10610 4375 10630 4395
rect 10655 4375 10675 4395
rect 10700 4375 10720 4395
<< metal1 >>
rect 295 6095 335 6500
rect 385 6475 425 6500
rect 385 6215 390 6475
rect 420 6215 425 6475
rect 295 6085 330 6095
rect 295 5815 300 6085
rect 295 5805 330 5815
rect -20 4905 275 4925
rect -20 4865 20 4905
rect 205 4400 245 4805
rect 205 4370 210 4400
rect 240 4370 245 4400
rect 205 1930 245 4370
rect 295 1930 335 5805
rect 385 1930 425 6215
rect 515 4905 11810 4925
rect 11770 4865 11810 4905
rect 1295 4410 1315 4415
rect 1835 4410 1855 4415
rect 2015 4410 2035 4415
rect 1110 4400 1140 4410
rect 1290 4400 1320 4410
rect 1830 4400 1860 4410
rect 2010 4400 2040 4410
rect 2510 4400 2530 4415
rect 2555 4410 2575 4415
rect 2640 4410 2670 4415
rect 2550 4400 2580 4410
rect 2645 4405 2665 4410
rect 2600 4400 2620 4405
rect 2690 4400 2710 4415
rect 2735 4410 2755 4415
rect 2730 4400 2760 4410
rect 2780 4400 2800 4405
rect 1270 4370 1275 4400
rect 1335 4370 1340 4400
rect 1810 4370 1815 4400
rect 1875 4370 1880 4400
rect 1990 4370 1995 4400
rect 2055 4370 2060 4400
rect 2510 4395 2535 4400
rect 2530 4375 2535 4395
rect 2510 4370 2535 4375
rect 2595 4395 2625 4400
rect 2595 4375 2600 4395
rect 2620 4375 2625 4395
rect 2595 4370 2625 4375
rect 2685 4395 2715 4400
rect 2685 4375 2690 4395
rect 2710 4375 2715 4395
rect 2685 4370 2715 4375
rect 2775 4395 2800 4400
rect 2775 4375 2780 4395
rect 2775 4370 2800 4375
rect 1110 4360 1140 4370
rect 1290 4360 1320 4370
rect 1830 4360 1860 4370
rect 2010 4360 2040 4370
rect 2510 4365 2530 4370
rect 2550 4360 2580 4370
rect 1295 4355 1315 4360
rect 1835 4355 1855 4360
rect 2015 4355 2035 4360
rect 2555 4355 2575 4360
rect 2600 4355 2620 4370
rect 2690 4365 2710 4370
rect 2730 4360 2760 4370
rect 2735 4355 2755 4360
rect 2780 4355 2800 4370
rect 3230 4400 3250 4415
rect 3275 4410 3295 4415
rect 3360 4410 3390 4415
rect 3270 4400 3300 4410
rect 3365 4405 3385 4410
rect 3320 4400 3340 4405
rect 3410 4400 3430 4415
rect 3455 4410 3475 4415
rect 3450 4400 3480 4410
rect 3500 4400 3520 4405
rect 3230 4395 3255 4400
rect 3250 4375 3255 4395
rect 3230 4370 3255 4375
rect 3315 4395 3345 4400
rect 3315 4375 3320 4395
rect 3340 4375 3345 4395
rect 3315 4370 3345 4375
rect 3405 4395 3435 4400
rect 3405 4375 3410 4395
rect 3430 4375 3435 4395
rect 3405 4370 3435 4375
rect 3495 4395 3520 4400
rect 3495 4375 3500 4395
rect 3495 4370 3520 4375
rect 3230 4365 3250 4370
rect 3270 4360 3300 4370
rect 3275 4355 3295 4360
rect 3320 4355 3340 4370
rect 3410 4365 3430 4370
rect 3450 4360 3480 4370
rect 3455 4355 3475 4360
rect 3500 4355 3520 4370
rect 3950 4400 3970 4415
rect 3995 4410 4015 4415
rect 4080 4410 4110 4415
rect 3990 4400 4020 4410
rect 4085 4405 4105 4410
rect 4040 4400 4060 4405
rect 4130 4400 4150 4415
rect 4175 4410 4195 4415
rect 4170 4400 4200 4410
rect 4220 4400 4240 4405
rect 3950 4395 3975 4400
rect 3970 4375 3975 4395
rect 3950 4370 3975 4375
rect 4035 4395 4065 4400
rect 4035 4375 4040 4395
rect 4060 4375 4065 4395
rect 4035 4370 4065 4375
rect 4125 4395 4155 4400
rect 4125 4375 4130 4395
rect 4150 4375 4155 4395
rect 4125 4370 4155 4375
rect 4215 4395 4240 4400
rect 4215 4375 4220 4395
rect 4215 4370 4240 4375
rect 3950 4365 3970 4370
rect 3990 4360 4020 4370
rect 3995 4355 4015 4360
rect 4040 4355 4060 4370
rect 4130 4365 4150 4370
rect 4170 4360 4200 4370
rect 4175 4355 4195 4360
rect 4220 4355 4240 4370
rect 7550 4400 7570 4415
rect 7595 4410 7615 4415
rect 7680 4410 7710 4415
rect 7590 4400 7620 4410
rect 7685 4405 7705 4410
rect 7640 4400 7660 4405
rect 7730 4400 7750 4415
rect 7775 4410 7795 4415
rect 7770 4400 7800 4410
rect 7820 4400 7840 4405
rect 7550 4395 7575 4400
rect 7570 4375 7575 4395
rect 7550 4370 7575 4375
rect 7635 4395 7665 4400
rect 7635 4375 7640 4395
rect 7660 4375 7665 4395
rect 7635 4370 7665 4375
rect 7725 4395 7755 4400
rect 7725 4375 7730 4395
rect 7750 4375 7755 4395
rect 7725 4370 7755 4375
rect 7815 4395 7840 4400
rect 7815 4375 7820 4395
rect 7815 4370 7840 4375
rect 7550 4365 7570 4370
rect 7590 4360 7620 4370
rect 7595 4355 7615 4360
rect 7640 4355 7660 4370
rect 7730 4365 7750 4370
rect 7770 4360 7800 4370
rect 7775 4355 7795 4360
rect 7820 4355 7840 4370
rect 8270 4400 8290 4415
rect 8315 4410 8335 4415
rect 8400 4410 8430 4415
rect 8310 4400 8340 4410
rect 8405 4405 8425 4410
rect 8360 4400 8380 4405
rect 8450 4400 8470 4415
rect 8495 4410 8515 4415
rect 8490 4400 8520 4410
rect 8540 4400 8560 4405
rect 8270 4395 8295 4400
rect 8290 4375 8295 4395
rect 8270 4370 8295 4375
rect 8355 4395 8385 4400
rect 8355 4375 8360 4395
rect 8380 4375 8385 4395
rect 8355 4370 8385 4375
rect 8445 4395 8475 4400
rect 8445 4375 8450 4395
rect 8470 4375 8475 4395
rect 8445 4370 8475 4375
rect 8535 4395 8560 4400
rect 8535 4375 8540 4395
rect 8535 4370 8560 4375
rect 8270 4365 8290 4370
rect 8310 4360 8340 4370
rect 8315 4355 8335 4360
rect 8360 4355 8380 4370
rect 8450 4365 8470 4370
rect 8490 4360 8520 4370
rect 8495 4355 8515 4360
rect 8540 4355 8560 4370
rect 8990 4400 9010 4415
rect 9035 4410 9055 4415
rect 9120 4410 9150 4415
rect 9030 4400 9060 4410
rect 9125 4405 9145 4410
rect 9080 4400 9100 4405
rect 9170 4400 9190 4415
rect 9215 4410 9235 4415
rect 9210 4400 9240 4410
rect 9260 4400 9280 4405
rect 8990 4395 9015 4400
rect 9010 4375 9015 4395
rect 8990 4370 9015 4375
rect 9075 4395 9105 4400
rect 9075 4375 9080 4395
rect 9100 4375 9105 4395
rect 9075 4370 9105 4375
rect 9165 4395 9195 4400
rect 9165 4375 9170 4395
rect 9190 4375 9195 4395
rect 9165 4370 9195 4375
rect 9255 4395 9280 4400
rect 9255 4375 9260 4395
rect 9255 4370 9280 4375
rect 8990 4365 9010 4370
rect 9030 4360 9060 4370
rect 9035 4355 9055 4360
rect 9080 4355 9100 4370
rect 9170 4365 9190 4370
rect 9210 4360 9240 4370
rect 9215 4355 9235 4360
rect 9260 4355 9280 4370
rect 9710 4400 9730 4415
rect 9755 4410 9775 4415
rect 9840 4410 9870 4415
rect 9750 4400 9780 4410
rect 9845 4405 9865 4410
rect 9800 4400 9820 4405
rect 9890 4400 9910 4415
rect 9935 4410 9955 4415
rect 9930 4400 9960 4410
rect 9980 4400 10000 4405
rect 9710 4395 9735 4400
rect 9730 4375 9735 4395
rect 9710 4370 9735 4375
rect 9795 4395 9825 4400
rect 9795 4375 9800 4395
rect 9820 4375 9825 4395
rect 9795 4370 9825 4375
rect 9885 4395 9915 4400
rect 9885 4375 9890 4395
rect 9910 4375 9915 4395
rect 9885 4370 9915 4375
rect 9975 4395 10000 4400
rect 9975 4375 9980 4395
rect 9975 4370 10000 4375
rect 9710 4365 9730 4370
rect 9750 4360 9780 4370
rect 9755 4355 9775 4360
rect 9800 4355 9820 4370
rect 9890 4365 9910 4370
rect 9930 4360 9960 4370
rect 9935 4355 9955 4360
rect 9980 4355 10000 4370
rect 10430 4400 10450 4415
rect 10475 4410 10495 4415
rect 10560 4410 10590 4415
rect 10470 4400 10500 4410
rect 10565 4405 10585 4410
rect 10520 4400 10540 4405
rect 10610 4400 10630 4415
rect 10655 4410 10675 4415
rect 10650 4400 10680 4410
rect 10700 4400 10720 4405
rect 10430 4395 10455 4400
rect 10450 4375 10455 4395
rect 10430 4370 10455 4375
rect 10515 4395 10545 4400
rect 10515 4375 10520 4395
rect 10540 4375 10545 4395
rect 10515 4370 10545 4375
rect 10605 4395 10635 4400
rect 10605 4375 10610 4395
rect 10630 4375 10635 4395
rect 10605 4370 10635 4375
rect 10695 4395 10720 4400
rect 10695 4375 10700 4395
rect 10695 4370 10720 4375
rect 10430 4365 10450 4370
rect 10470 4360 10500 4370
rect 10475 4355 10495 4360
rect 10520 4355 10540 4370
rect 10610 4365 10630 4370
rect 10650 4360 10680 4370
rect 10655 4355 10675 4360
rect 10700 4355 10720 4370
rect 11285 605 11305 4865
rect 11375 605 11395 4865
rect 11465 605 11485 4865
rect 11555 605 11575 4865
<< via1 >>
rect 390 6470 420 6475
rect 390 6220 395 6470
rect 395 6220 415 6470
rect 415 6220 420 6470
rect 390 6215 420 6220
rect 300 6080 330 6085
rect 300 5820 305 6080
rect 305 5820 325 6080
rect 325 5820 330 6080
rect 300 5815 330 5820
rect 210 4370 240 4400
rect 1110 4370 1140 4400
rect 1290 4395 1320 4400
rect 1290 4375 1295 4395
rect 1295 4375 1315 4395
rect 1315 4375 1320 4395
rect 1290 4370 1320 4375
rect 1830 4395 1860 4400
rect 1830 4375 1835 4395
rect 1835 4375 1855 4395
rect 1855 4375 1860 4395
rect 1830 4370 1860 4375
rect 2010 4395 2040 4400
rect 2010 4375 2015 4395
rect 2015 4375 2035 4395
rect 2035 4375 2040 4395
rect 2010 4370 2040 4375
rect 2550 4395 2580 4400
rect 2550 4375 2555 4395
rect 2555 4375 2575 4395
rect 2575 4375 2580 4395
rect 2550 4370 2580 4375
rect 2730 4395 2760 4400
rect 2730 4375 2735 4395
rect 2735 4375 2755 4395
rect 2755 4375 2760 4395
rect 2730 4370 2760 4375
rect 3270 4395 3300 4400
rect 3270 4375 3275 4395
rect 3275 4375 3295 4395
rect 3295 4375 3300 4395
rect 3270 4370 3300 4375
rect 3450 4395 3480 4400
rect 3450 4375 3455 4395
rect 3455 4375 3475 4395
rect 3475 4375 3480 4395
rect 3450 4370 3480 4375
rect 3990 4395 4020 4400
rect 3990 4375 3995 4395
rect 3995 4375 4015 4395
rect 4015 4375 4020 4395
rect 3990 4370 4020 4375
rect 4170 4395 4200 4400
rect 4170 4375 4175 4395
rect 4175 4375 4195 4395
rect 4195 4375 4200 4395
rect 4170 4370 4200 4375
rect 7590 4395 7620 4400
rect 7590 4375 7595 4395
rect 7595 4375 7615 4395
rect 7615 4375 7620 4395
rect 7590 4370 7620 4375
rect 7770 4395 7800 4400
rect 7770 4375 7775 4395
rect 7775 4375 7795 4395
rect 7795 4375 7800 4395
rect 7770 4370 7800 4375
rect 8310 4395 8340 4400
rect 8310 4375 8315 4395
rect 8315 4375 8335 4395
rect 8335 4375 8340 4395
rect 8310 4370 8340 4375
rect 8490 4395 8520 4400
rect 8490 4375 8495 4395
rect 8495 4375 8515 4395
rect 8515 4375 8520 4395
rect 8490 4370 8520 4375
rect 9030 4395 9060 4400
rect 9030 4375 9035 4395
rect 9035 4375 9055 4395
rect 9055 4375 9060 4395
rect 9030 4370 9060 4375
rect 9210 4395 9240 4400
rect 9210 4375 9215 4395
rect 9215 4375 9235 4395
rect 9235 4375 9240 4395
rect 9210 4370 9240 4375
rect 9750 4395 9780 4400
rect 9750 4375 9755 4395
rect 9755 4375 9775 4395
rect 9775 4375 9780 4395
rect 9750 4370 9780 4375
rect 9930 4395 9960 4400
rect 9930 4375 9935 4395
rect 9935 4375 9955 4395
rect 9955 4375 9960 4395
rect 9930 4370 9960 4375
rect 10470 4395 10500 4400
rect 10470 4375 10475 4395
rect 10475 4375 10495 4395
rect 10495 4375 10500 4395
rect 10470 4370 10500 4375
rect 10650 4395 10680 4400
rect 10650 4375 10655 4395
rect 10655 4375 10675 4395
rect 10675 4375 10680 4395
rect 10650 4370 10680 4375
<< metal2 >>
rect 380 6485 430 6490
rect 380 6205 385 6485
rect 425 6205 430 6485
rect 380 6200 430 6205
rect 290 6095 340 6100
rect 290 5805 295 6095
rect 335 5805 340 6095
rect 290 5800 340 5805
rect 145 4925 665 4930
rect -800 4915 12600 4925
rect -800 4835 -790 4915
rect -510 4835 12310 4915
rect 12590 4835 12600 4915
rect -800 4825 12600 4835
rect 115 4410 11675 4415
rect 115 4400 1105 4410
rect 115 4370 210 4400
rect 240 4370 1105 4400
rect 115 4360 1105 4370
rect 1145 4360 1285 4410
rect 1325 4360 1825 4410
rect 1865 4360 2005 4410
rect 2045 4360 2545 4410
rect 2585 4360 2725 4410
rect 2765 4360 3265 4410
rect 3305 4360 3445 4410
rect 3485 4360 3985 4410
rect 4025 4360 4165 4410
rect 4205 4360 7585 4410
rect 7625 4360 7765 4410
rect 7805 4360 8305 4410
rect 8345 4360 8485 4410
rect 8525 4360 9025 4410
rect 9065 4360 9205 4410
rect 9245 4360 9745 4410
rect 9785 4360 9925 4410
rect 9965 4360 10465 4410
rect 10505 4360 10645 4410
rect 10685 4360 11675 4410
rect 115 4355 11675 4360
rect -800 3935 12600 3945
rect -800 3855 -390 3935
rect -110 3855 11910 3935
rect 12190 3855 12600 3935
rect -800 3845 12600 3855
rect -800 2920 12600 2930
rect -800 2840 -790 2920
rect -510 2840 12310 2920
rect 12590 2840 12600 2920
rect -800 2830 12600 2840
rect -800 1900 12600 1910
rect -800 1820 -390 1900
rect -110 1820 11910 1900
rect 12190 1820 12600 1900
rect -800 1810 12600 1820
rect -800 960 12600 970
rect -800 880 -790 960
rect -510 880 12310 960
rect 12590 880 12600 960
rect -800 870 12600 880
rect -800 20 12600 30
rect -800 -60 -390 20
rect -110 -60 11910 20
rect 12190 -60 12600 20
rect -800 -70 12600 -60
<< via2 >>
rect 385 6475 425 6485
rect 385 6215 390 6475
rect 390 6215 420 6475
rect 420 6215 425 6475
rect 385 6205 425 6215
rect 295 6085 335 6095
rect 295 5815 300 6085
rect 300 5815 330 6085
rect 330 5815 335 6085
rect 295 5805 335 5815
rect -790 4835 -510 4915
rect 12310 4835 12590 4915
rect 1105 4400 1145 4410
rect 1105 4370 1110 4400
rect 1110 4370 1140 4400
rect 1140 4370 1145 4400
rect 1105 4360 1145 4370
rect 1285 4400 1325 4410
rect 1285 4370 1290 4400
rect 1290 4370 1320 4400
rect 1320 4370 1325 4400
rect 1285 4360 1325 4370
rect 1825 4400 1865 4410
rect 1825 4370 1830 4400
rect 1830 4370 1860 4400
rect 1860 4370 1865 4400
rect 1825 4360 1865 4370
rect 2005 4400 2045 4410
rect 2005 4370 2010 4400
rect 2010 4370 2040 4400
rect 2040 4370 2045 4400
rect 2005 4360 2045 4370
rect 2545 4400 2585 4410
rect 2545 4370 2550 4400
rect 2550 4370 2580 4400
rect 2580 4370 2585 4400
rect 2545 4360 2585 4370
rect 2725 4400 2765 4410
rect 2725 4370 2730 4400
rect 2730 4370 2760 4400
rect 2760 4370 2765 4400
rect 2725 4360 2765 4370
rect 3265 4400 3305 4410
rect 3265 4370 3270 4400
rect 3270 4370 3300 4400
rect 3300 4370 3305 4400
rect 3265 4360 3305 4370
rect 3445 4400 3485 4410
rect 3445 4370 3450 4400
rect 3450 4370 3480 4400
rect 3480 4370 3485 4400
rect 3445 4360 3485 4370
rect 3985 4400 4025 4410
rect 3985 4370 3990 4400
rect 3990 4370 4020 4400
rect 4020 4370 4025 4400
rect 3985 4360 4025 4370
rect 4165 4400 4205 4410
rect 4165 4370 4170 4400
rect 4170 4370 4200 4400
rect 4200 4370 4205 4400
rect 4165 4360 4205 4370
rect 7585 4400 7625 4410
rect 7585 4370 7590 4400
rect 7590 4370 7620 4400
rect 7620 4370 7625 4400
rect 7585 4360 7625 4370
rect 7765 4400 7805 4410
rect 7765 4370 7770 4400
rect 7770 4370 7800 4400
rect 7800 4370 7805 4400
rect 7765 4360 7805 4370
rect 8305 4400 8345 4410
rect 8305 4370 8310 4400
rect 8310 4370 8340 4400
rect 8340 4370 8345 4400
rect 8305 4360 8345 4370
rect 8485 4400 8525 4410
rect 8485 4370 8490 4400
rect 8490 4370 8520 4400
rect 8520 4370 8525 4400
rect 8485 4360 8525 4370
rect 9025 4400 9065 4410
rect 9025 4370 9030 4400
rect 9030 4370 9060 4400
rect 9060 4370 9065 4400
rect 9025 4360 9065 4370
rect 9205 4400 9245 4410
rect 9205 4370 9210 4400
rect 9210 4370 9240 4400
rect 9240 4370 9245 4400
rect 9205 4360 9245 4370
rect 9745 4400 9785 4410
rect 9745 4370 9750 4400
rect 9750 4370 9780 4400
rect 9780 4370 9785 4400
rect 9745 4360 9785 4370
rect 9925 4400 9965 4410
rect 9925 4370 9930 4400
rect 9930 4370 9960 4400
rect 9960 4370 9965 4400
rect 9925 4360 9965 4370
rect 10465 4400 10505 4410
rect 10465 4370 10470 4400
rect 10470 4370 10500 4400
rect 10500 4370 10505 4400
rect 10465 4360 10505 4370
rect 10645 4400 10685 4410
rect 10645 4370 10650 4400
rect 10650 4370 10680 4400
rect 10680 4370 10685 4400
rect 10645 4360 10685 4370
rect -390 3855 -110 3935
rect 11910 3855 12190 3935
rect -790 2840 -510 2920
rect 12310 2840 12590 2920
rect -390 1820 -110 1900
rect 11910 1820 12190 1900
rect -790 880 -510 960
rect 12310 880 12590 960
rect -390 -60 -110 20
rect 11910 -60 12190 20
<< metal3 >>
rect 380 6485 430 6490
rect 380 6205 385 6485
rect 425 6205 430 6485
rect 380 6200 430 6205
rect 290 6095 340 6100
rect 290 5805 295 6095
rect 335 5805 340 6095
rect 290 5800 340 5805
rect -800 5650 -500 5700
rect -800 5450 -750 5650
rect -550 5450 -500 5650
rect -800 4915 -500 5450
rect -800 4835 -790 4915
rect -510 4835 -500 4915
rect -800 2920 -500 4835
rect -800 2840 -790 2920
rect -510 2840 -500 2920
rect -800 960 -500 2840
rect -800 880 -790 960
rect -510 880 -500 960
rect -800 -650 -500 880
rect -800 -850 -750 -650
rect -550 -850 -500 -650
rect -800 -900 -500 -850
rect -400 5250 -100 5300
rect -400 5050 -350 5250
rect -150 5050 -100 5250
rect -400 3935 -100 5050
rect 11900 5250 12200 6500
rect 11900 5050 11950 5250
rect 12150 5050 12200 5250
rect 1100 4410 1150 4415
rect 1100 4360 1105 4410
rect 1145 4360 1150 4410
rect 1100 4355 1150 4360
rect 1280 4410 1330 4415
rect 1280 4360 1285 4410
rect 1325 4360 1330 4410
rect 1280 4355 1330 4360
rect 1820 4410 1870 4415
rect 1820 4360 1825 4410
rect 1865 4360 1870 4410
rect 1820 4355 1870 4360
rect 2000 4410 2050 4415
rect 2000 4360 2005 4410
rect 2045 4360 2050 4410
rect 2000 4355 2050 4360
rect 2540 4410 2590 4415
rect 2540 4360 2545 4410
rect 2585 4360 2590 4410
rect 2540 4355 2590 4360
rect 2720 4410 2770 4415
rect 2720 4360 2725 4410
rect 2765 4360 2770 4410
rect 2720 4355 2770 4360
rect 3260 4410 3310 4415
rect 3260 4360 3265 4410
rect 3305 4360 3310 4410
rect 3260 4355 3310 4360
rect 3440 4410 3490 4415
rect 3440 4360 3445 4410
rect 3485 4360 3490 4410
rect 3440 4355 3490 4360
rect 3980 4410 4030 4415
rect 3980 4360 3985 4410
rect 4025 4360 4030 4410
rect 3980 4355 4030 4360
rect 4160 4410 4210 4415
rect 4160 4360 4165 4410
rect 4205 4360 4210 4410
rect 4160 4355 4210 4360
rect 7580 4410 7630 4415
rect 7580 4360 7585 4410
rect 7625 4360 7630 4410
rect 7580 4355 7630 4360
rect 7760 4410 7810 4415
rect 7760 4360 7765 4410
rect 7805 4360 7810 4410
rect 7760 4355 7810 4360
rect 8300 4410 8350 4415
rect 8300 4360 8305 4410
rect 8345 4360 8350 4410
rect 8300 4355 8350 4360
rect 8480 4410 8530 4415
rect 8480 4360 8485 4410
rect 8525 4360 8530 4410
rect 8480 4355 8530 4360
rect 9020 4410 9070 4415
rect 9020 4360 9025 4410
rect 9065 4360 9070 4410
rect 9020 4355 9070 4360
rect 9200 4410 9250 4415
rect 9200 4360 9205 4410
rect 9245 4360 9250 4410
rect 9200 4355 9250 4360
rect 9740 4410 9790 4415
rect 9740 4360 9745 4410
rect 9785 4360 9790 4410
rect 9740 4355 9790 4360
rect 9920 4410 9970 4415
rect 9920 4360 9925 4410
rect 9965 4360 9970 4410
rect 9920 4355 9970 4360
rect 10460 4410 10510 4415
rect 10460 4360 10465 4410
rect 10505 4360 10510 4410
rect 10460 4355 10510 4360
rect 10640 4410 10690 4415
rect 10640 4360 10645 4410
rect 10685 4360 10690 4410
rect 10640 4355 10690 4360
rect -400 3855 -390 3935
rect -110 3855 -100 3935
rect -400 1900 -100 3855
rect -400 1820 -390 1900
rect -110 1820 -100 1900
rect -400 20 -100 1820
rect -400 -60 -390 20
rect -110 -60 -100 20
rect -400 -250 -100 -60
rect -400 -450 -350 -250
rect -150 -450 -100 -250
rect -400 -900 -100 -450
rect 11900 3935 12200 5050
rect 11900 3855 11910 3935
rect 12190 3855 12200 3935
rect 11900 1900 12200 3855
rect 11900 1820 11910 1900
rect 12190 1820 12200 1900
rect 11900 20 12200 1820
rect 11900 -60 11910 20
rect 12190 -60 12200 20
rect 11900 -250 12200 -60
rect 11900 -450 11950 -250
rect 12150 -450 12200 -250
rect 11900 -900 12200 -450
rect 12300 5650 12600 6500
rect 12300 5450 12350 5650
rect 12550 5450 12600 5650
rect 12300 4915 12600 5450
rect 12300 4835 12310 4915
rect 12590 4835 12600 4915
rect 12300 2920 12600 4835
rect 12300 2840 12310 2920
rect 12590 2840 12600 2920
rect 12300 960 12600 2840
rect 12300 880 12310 960
rect 12590 880 12600 960
rect 12300 -650 12600 880
rect 12300 -850 12350 -650
rect 12550 -850 12600 -650
rect 12300 -900 12600 -850
rect 12700 4450 13000 6500
rect 12700 4250 12750 4450
rect 12950 4250 13000 4450
rect 12700 -900 13000 4250
rect 13100 -900 13400 6500
rect 13500 -900 13800 6500
<< via3 >>
rect 385 6205 425 6485
rect 295 5805 335 6095
rect -750 5450 -550 5650
rect -750 -850 -550 -650
rect -350 5050 -150 5250
rect 11950 5050 12150 5250
rect -350 -450 -150 -250
rect 11950 -450 12150 -250
rect 12350 5450 12550 5650
rect 12350 -850 12550 -650
rect 12750 4250 12950 4450
<< metal4 >>
rect -800 6485 14100 6500
rect -800 6205 385 6485
rect 425 6205 14100 6485
rect -800 6200 14100 6205
rect -800 6095 14100 6100
rect -800 5805 295 6095
rect 335 5805 14100 6095
rect -800 5800 14100 5805
rect -800 5650 14100 5700
rect -800 5450 -750 5650
rect -550 5450 12350 5650
rect 12550 5450 14100 5650
rect -800 5400 14100 5450
rect -800 5250 14100 5300
rect -800 5050 -350 5250
rect -150 5050 11950 5250
rect 12150 5050 14100 5250
rect -800 5000 14100 5050
rect -800 4450 14100 4500
rect -800 4250 12750 4450
rect 12950 4250 14100 4450
rect -800 4200 14100 4250
rect -245 4195 715 4200
rect -800 -250 12600 -200
rect -800 -450 -350 -250
rect -150 -450 11950 -250
rect 12150 -450 12600 -250
rect -800 -500 12600 -450
rect -800 -650 12600 -600
rect -800 -850 -750 -650
rect -550 -850 12350 -650
rect 12550 -850 12600 -650
rect -800 -900 12600 -850
use buffer  buffer_0
timestamp 1624076896
transform 1 0 -9060 0 1 490
box 9040 3415 20870 4385
use ota  ota_0
timestamp 1624070110
transform 1 0 11680 0 1 1880
box -11700 -10 130 2005
use bias  bias_0
timestamp 1624062196
transform 1 0 465 0 1 0
box -485 -10 11350 1850
<< labels >>
rlabel metal4 14000 5400 14100 5700 1 VDDA
port 1 n
rlabel metal4 14000 5000 14100 5300 1 VSSA
port 2 n
rlabel metal4 14000 5800 14100 6100 1 INM
port 3 n
rlabel metal4 14000 6200 14100 6500 1 INP
port 4 n
rlabel metal4 14000 4200 14100 4500 1 OUT
port 5 n
rlabel metal1 225 4525 225 4525 1 X
rlabel metal1 11295 1310 11295 1310 1 P1
rlabel metal1 11385 1310 11385 1310 1 P2
rlabel metal1 11475 1310 11475 1310 1 N2
rlabel metal1 11565 1310 11565 1310 1 N1
<< end >>
