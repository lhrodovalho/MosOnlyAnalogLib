magic
tech sky130A
timestamp 1624051598
<< nwell >>
rect 10345 4105 12840 4385
<< mvnmos >>
rect 10455 3475 10505 3575
rect 10545 3475 10595 3575
rect 10635 3475 10685 3575
rect 10725 3475 10775 3575
rect 10815 3475 10865 3575
rect 10905 3475 10955 3575
rect 10995 3475 11045 3575
rect 11085 3475 11135 3575
rect 11175 3475 11225 3575
rect 11265 3475 11315 3575
rect 11355 3475 11405 3575
rect 11445 3475 11495 3575
rect 11535 3475 11585 3575
rect 11625 3475 11675 3575
rect 11715 3475 11765 3575
rect 11805 3475 11855 3575
rect 11895 3475 11945 3575
rect 11985 3475 12035 3575
rect 12075 3475 12125 3575
rect 12165 3475 12215 3575
rect 12255 3475 12305 3575
rect 12345 3475 12395 3575
rect 12435 3475 12485 3575
rect 12525 3475 12575 3575
rect 12615 3475 12665 3575
rect 12705 3475 12755 3575
<< mvpmos >>
rect 10455 4215 10505 4315
rect 10545 4215 10595 4315
rect 10635 4215 10685 4315
rect 10725 4215 10775 4315
rect 10815 4215 10865 4315
rect 10905 4215 10955 4315
rect 10995 4215 11045 4315
rect 11085 4215 11135 4315
rect 11175 4215 11225 4315
rect 11265 4215 11315 4315
rect 11355 4215 11405 4315
rect 11445 4215 11495 4315
rect 11535 4215 11585 4315
rect 11625 4215 11675 4315
rect 11715 4215 11765 4315
rect 11805 4215 11855 4315
rect 11895 4215 11945 4315
rect 11985 4215 12035 4315
rect 12075 4215 12125 4315
rect 12165 4215 12215 4315
rect 12255 4215 12305 4315
rect 12345 4215 12395 4315
rect 12435 4215 12485 4315
rect 12525 4215 12575 4315
rect 12615 4215 12665 4315
rect 12705 4215 12755 4315
<< mvndiff >>
rect 10415 3565 10455 3575
rect 10415 3485 10425 3565
rect 10445 3485 10455 3565
rect 10415 3475 10455 3485
rect 10505 3565 10545 3575
rect 10505 3485 10515 3565
rect 10535 3485 10545 3565
rect 10505 3475 10545 3485
rect 10595 3565 10635 3575
rect 10595 3485 10605 3565
rect 10625 3485 10635 3565
rect 10595 3475 10635 3485
rect 10685 3565 10725 3575
rect 10685 3485 10695 3565
rect 10715 3485 10725 3565
rect 10685 3475 10725 3485
rect 10775 3565 10815 3575
rect 10775 3485 10785 3565
rect 10805 3485 10815 3565
rect 10775 3475 10815 3485
rect 10865 3565 10905 3575
rect 10865 3485 10875 3565
rect 10895 3485 10905 3565
rect 10865 3475 10905 3485
rect 10955 3565 10995 3575
rect 10955 3485 10965 3565
rect 10985 3485 10995 3565
rect 10955 3475 10995 3485
rect 11045 3565 11085 3575
rect 11045 3485 11055 3565
rect 11075 3485 11085 3565
rect 11045 3475 11085 3485
rect 11135 3565 11175 3575
rect 11135 3485 11145 3565
rect 11165 3485 11175 3565
rect 11135 3475 11175 3485
rect 11225 3565 11265 3575
rect 11225 3485 11235 3565
rect 11255 3485 11265 3565
rect 11225 3475 11265 3485
rect 11315 3565 11355 3575
rect 11315 3485 11325 3565
rect 11345 3485 11355 3565
rect 11315 3475 11355 3485
rect 11405 3565 11445 3575
rect 11405 3485 11415 3565
rect 11435 3485 11445 3565
rect 11405 3475 11445 3485
rect 11495 3565 11535 3575
rect 11495 3485 11505 3565
rect 11525 3485 11535 3565
rect 11495 3475 11535 3485
rect 11585 3565 11625 3575
rect 11585 3485 11595 3565
rect 11615 3485 11625 3565
rect 11585 3475 11625 3485
rect 11675 3565 11715 3575
rect 11675 3485 11685 3565
rect 11705 3485 11715 3565
rect 11675 3475 11715 3485
rect 11765 3565 11805 3575
rect 11765 3485 11775 3565
rect 11795 3485 11805 3565
rect 11765 3475 11805 3485
rect 11855 3565 11895 3575
rect 11855 3485 11865 3565
rect 11885 3485 11895 3565
rect 11855 3475 11895 3485
rect 11945 3565 11985 3575
rect 11945 3485 11955 3565
rect 11975 3485 11985 3565
rect 11945 3475 11985 3485
rect 12035 3565 12075 3575
rect 12035 3485 12045 3565
rect 12065 3485 12075 3565
rect 12035 3475 12075 3485
rect 12125 3565 12165 3575
rect 12125 3485 12135 3565
rect 12155 3485 12165 3565
rect 12125 3475 12165 3485
rect 12215 3565 12255 3575
rect 12215 3485 12225 3565
rect 12245 3485 12255 3565
rect 12215 3475 12255 3485
rect 12305 3565 12345 3575
rect 12305 3485 12315 3565
rect 12335 3485 12345 3565
rect 12305 3475 12345 3485
rect 12395 3565 12435 3575
rect 12395 3485 12405 3565
rect 12425 3485 12435 3565
rect 12395 3475 12435 3485
rect 12485 3565 12525 3575
rect 12485 3485 12495 3565
rect 12515 3485 12525 3565
rect 12485 3475 12525 3485
rect 12575 3565 12615 3575
rect 12575 3485 12585 3565
rect 12605 3485 12615 3565
rect 12575 3475 12615 3485
rect 12665 3565 12705 3575
rect 12665 3485 12675 3565
rect 12695 3485 12705 3565
rect 12665 3475 12705 3485
rect 12755 3565 12794 3575
rect 12755 3485 12765 3565
rect 12785 3485 12794 3565
rect 12755 3475 12794 3485
<< mvpdiff >>
rect 10415 4305 10455 4315
rect 10415 4225 10425 4305
rect 10445 4225 10455 4305
rect 10415 4215 10455 4225
rect 10505 4305 10545 4315
rect 10505 4225 10515 4305
rect 10535 4225 10545 4305
rect 10505 4215 10545 4225
rect 10595 4305 10635 4315
rect 10595 4225 10605 4305
rect 10625 4225 10635 4305
rect 10595 4215 10635 4225
rect 10685 4305 10725 4315
rect 10685 4225 10695 4305
rect 10715 4225 10725 4305
rect 10685 4215 10725 4225
rect 10775 4305 10815 4315
rect 10775 4225 10785 4305
rect 10805 4225 10815 4305
rect 10775 4215 10815 4225
rect 10865 4305 10905 4315
rect 10865 4225 10875 4305
rect 10895 4225 10905 4305
rect 10865 4215 10905 4225
rect 10955 4305 10995 4315
rect 10955 4225 10965 4305
rect 10985 4225 10995 4305
rect 10955 4215 10995 4225
rect 11045 4305 11085 4315
rect 11045 4225 11055 4305
rect 11075 4225 11085 4305
rect 11045 4215 11085 4225
rect 11135 4305 11175 4315
rect 11135 4225 11145 4305
rect 11165 4225 11175 4305
rect 11135 4215 11175 4225
rect 11225 4305 11265 4315
rect 11225 4225 11235 4305
rect 11255 4225 11265 4305
rect 11225 4215 11265 4225
rect 11315 4305 11355 4315
rect 11315 4225 11325 4305
rect 11345 4225 11355 4305
rect 11315 4215 11355 4225
rect 11405 4305 11445 4315
rect 11405 4225 11415 4305
rect 11435 4225 11445 4305
rect 11405 4215 11445 4225
rect 11495 4305 11535 4315
rect 11495 4225 11505 4305
rect 11525 4225 11535 4305
rect 11495 4215 11535 4225
rect 11585 4305 11625 4315
rect 11585 4225 11595 4305
rect 11615 4225 11625 4305
rect 11585 4215 11625 4225
rect 11675 4305 11715 4315
rect 11675 4225 11685 4305
rect 11705 4225 11715 4305
rect 11675 4215 11715 4225
rect 11765 4305 11805 4315
rect 11765 4225 11775 4305
rect 11795 4225 11805 4305
rect 11765 4215 11805 4225
rect 11855 4305 11895 4315
rect 11855 4225 11865 4305
rect 11885 4225 11895 4305
rect 11855 4215 11895 4225
rect 11945 4305 11985 4315
rect 11945 4225 11955 4305
rect 11975 4225 11985 4305
rect 11945 4215 11985 4225
rect 12035 4305 12075 4315
rect 12035 4225 12045 4305
rect 12065 4225 12075 4305
rect 12035 4215 12075 4225
rect 12125 4305 12165 4315
rect 12125 4225 12135 4305
rect 12155 4225 12165 4305
rect 12125 4215 12165 4225
rect 12215 4305 12255 4315
rect 12215 4225 12225 4305
rect 12245 4225 12255 4305
rect 12215 4215 12255 4225
rect 12305 4305 12345 4315
rect 12305 4225 12315 4305
rect 12335 4225 12345 4305
rect 12305 4215 12345 4225
rect 12395 4305 12435 4315
rect 12395 4225 12405 4305
rect 12425 4225 12435 4305
rect 12395 4215 12435 4225
rect 12485 4305 12525 4315
rect 12485 4225 12495 4305
rect 12515 4225 12525 4305
rect 12485 4215 12525 4225
rect 12575 4305 12615 4315
rect 12575 4225 12585 4305
rect 12605 4225 12615 4305
rect 12575 4215 12615 4225
rect 12665 4305 12705 4315
rect 12665 4225 12675 4305
rect 12695 4225 12705 4305
rect 12665 4215 12705 4225
rect 12755 4305 12794 4315
rect 12755 4225 12765 4305
rect 12785 4225 12794 4305
rect 12755 4215 12794 4225
<< mvndiffc >>
rect 10425 3485 10445 3565
rect 10515 3485 10535 3565
rect 10605 3485 10625 3565
rect 10695 3485 10715 3565
rect 10785 3485 10805 3565
rect 10875 3485 10895 3565
rect 10965 3485 10985 3565
rect 11055 3485 11075 3565
rect 11145 3485 11165 3565
rect 11235 3485 11255 3565
rect 11325 3485 11345 3565
rect 11415 3485 11435 3565
rect 11505 3485 11525 3565
rect 11595 3485 11615 3565
rect 11685 3485 11705 3565
rect 11775 3485 11795 3565
rect 11865 3485 11885 3565
rect 11955 3485 11975 3565
rect 12045 3485 12065 3565
rect 12135 3485 12155 3565
rect 12225 3485 12245 3565
rect 12315 3485 12335 3565
rect 12405 3485 12425 3565
rect 12495 3485 12515 3565
rect 12585 3485 12605 3565
rect 12675 3485 12695 3565
rect 12765 3485 12785 3565
<< mvpdiffc >>
rect 10425 4225 10445 4305
rect 10515 4225 10535 4305
rect 10605 4225 10625 4305
rect 10695 4225 10715 4305
rect 10785 4225 10805 4305
rect 10875 4225 10895 4305
rect 10965 4225 10985 4305
rect 11055 4225 11075 4305
rect 11145 4225 11165 4305
rect 11235 4225 11255 4305
rect 11325 4225 11345 4305
rect 11415 4225 11435 4305
rect 11505 4225 11525 4305
rect 11595 4225 11615 4305
rect 11685 4225 11705 4305
rect 11775 4225 11795 4305
rect 11865 4225 11885 4305
rect 11955 4225 11975 4305
rect 12045 4225 12065 4305
rect 12135 4225 12155 4305
rect 12225 4225 12245 4305
rect 12315 4225 12335 4305
rect 12405 4225 12425 4305
rect 12495 4225 12515 4305
rect 12585 4225 12605 4305
rect 12675 4225 12695 4305
rect 12765 4225 12785 4305
<< psubdiff >>
rect 10290 4065 10310 4375
rect 10290 4045 10470 4065
rect 10490 4045 10560 4065
rect 10580 4045 10650 4065
rect 10670 4045 10740 4065
rect 10760 4045 10830 4065
rect 10850 4045 10920 4065
rect 10940 4045 11010 4065
rect 11030 4045 11100 4065
rect 11120 4045 11190 4065
rect 11210 4045 11280 4065
rect 11300 4045 11370 4065
rect 11390 4045 11460 4065
rect 11480 4045 11550 4065
rect 11570 4045 11640 4065
rect 11660 4045 11730 4065
rect 11750 4045 11820 4065
rect 11840 4045 11910 4065
rect 11930 4045 12000 4065
rect 12020 4045 12090 4065
rect 12110 4045 12180 4065
rect 12200 4045 12270 4065
rect 12290 4045 12360 4065
rect 12380 4045 12450 4065
rect 12470 4045 12540 4065
rect 12560 4045 12630 4065
rect 12650 4045 12720 4065
rect 12740 4045 12794 4065
rect 10290 3645 10470 3665
rect 10490 3645 10560 3665
rect 10580 3645 10650 3665
rect 10670 3645 10740 3665
rect 10760 3645 10830 3665
rect 10850 3645 10920 3665
rect 10940 3645 11010 3665
rect 11030 3645 11100 3665
rect 11120 3645 11190 3665
rect 11210 3645 11280 3665
rect 11300 3645 11370 3665
rect 11390 3645 11460 3665
rect 11480 3645 11550 3665
rect 11570 3645 11640 3665
rect 11660 3645 11730 3665
rect 11750 3645 11820 3665
rect 11840 3645 11910 3665
rect 11930 3645 12000 3665
rect 12020 3645 12090 3665
rect 12110 3645 12180 3665
rect 12200 3645 12270 3665
rect 12290 3645 12360 3665
rect 12380 3645 12450 3665
rect 12470 3645 12540 3665
rect 12560 3645 12630 3665
rect 12650 3645 12720 3665
rect 12740 3645 12794 3665
rect 10290 3445 10310 3645
rect 10280 3425 10470 3445
rect 10490 3425 10560 3445
rect 10580 3425 10650 3445
rect 10670 3425 10740 3445
rect 10760 3425 10830 3445
rect 10850 3425 10920 3445
rect 10940 3425 11010 3445
rect 11030 3425 11100 3445
rect 11120 3425 11190 3445
rect 11210 3425 11280 3445
rect 11300 3425 11370 3445
rect 11390 3425 11460 3445
rect 11480 3425 11550 3445
rect 11570 3425 11640 3445
rect 11660 3425 11730 3445
rect 11750 3425 11820 3445
rect 11840 3425 11910 3445
rect 11930 3425 12000 3445
rect 12020 3425 12090 3445
rect 12110 3425 12180 3445
rect 12200 3425 12270 3445
rect 12290 3425 12360 3445
rect 12380 3425 12450 3445
rect 12470 3425 12540 3445
rect 12560 3425 12630 3445
rect 12650 3425 12720 3445
rect 12740 3425 12794 3445
<< nsubdiff >>
rect 10365 4345 10470 4365
rect 10490 4345 10560 4365
rect 10580 4345 10650 4365
rect 10670 4345 10740 4365
rect 10760 4345 10830 4365
rect 10850 4345 10920 4365
rect 10940 4345 11010 4365
rect 11030 4345 11100 4365
rect 11120 4345 11190 4365
rect 11210 4345 11280 4365
rect 11300 4345 11370 4365
rect 11390 4345 11460 4365
rect 11480 4345 11550 4365
rect 11570 4345 11640 4365
rect 11660 4345 11730 4365
rect 11750 4345 11820 4365
rect 11840 4345 11910 4365
rect 11930 4345 12000 4365
rect 12020 4345 12090 4365
rect 12110 4345 12180 4365
rect 12200 4345 12270 4365
rect 12290 4345 12360 4365
rect 12380 4345 12450 4365
rect 12470 4345 12540 4365
rect 12560 4345 12630 4365
rect 12650 4345 12720 4365
rect 12740 4345 12794 4365
rect 10365 4145 10385 4345
rect 10365 4125 10470 4145
rect 10490 4125 10560 4145
rect 10580 4125 10650 4145
rect 10670 4125 10740 4145
rect 10760 4125 10830 4145
rect 10850 4125 10920 4145
rect 10940 4125 11010 4145
rect 11030 4125 11100 4145
rect 11120 4125 11190 4145
rect 11210 4125 11280 4145
rect 11300 4125 11370 4145
rect 11390 4125 11460 4145
rect 11480 4125 11550 4145
rect 11570 4125 11640 4145
rect 11660 4125 11730 4145
rect 11750 4125 11820 4145
rect 11840 4125 11910 4145
rect 11930 4125 12000 4145
rect 12020 4125 12090 4145
rect 12110 4125 12180 4145
rect 12200 4125 12270 4145
rect 12290 4125 12360 4145
rect 12380 4125 12450 4145
rect 12470 4125 12540 4145
rect 12560 4125 12630 4145
rect 12650 4125 12720 4145
rect 12740 4125 12794 4145
<< psubdiffcont >>
rect 10470 4045 10490 4065
rect 10560 4045 10580 4065
rect 10650 4045 10670 4065
rect 10740 4045 10760 4065
rect 10830 4045 10850 4065
rect 10920 4045 10940 4065
rect 11010 4045 11030 4065
rect 11100 4045 11120 4065
rect 11190 4045 11210 4065
rect 11280 4045 11300 4065
rect 11370 4045 11390 4065
rect 11460 4045 11480 4065
rect 11550 4045 11570 4065
rect 11640 4045 11660 4065
rect 11730 4045 11750 4065
rect 11820 4045 11840 4065
rect 11910 4045 11930 4065
rect 12000 4045 12020 4065
rect 12090 4045 12110 4065
rect 12180 4045 12200 4065
rect 12270 4045 12290 4065
rect 12360 4045 12380 4065
rect 12450 4045 12470 4065
rect 12540 4045 12560 4065
rect 12630 4045 12650 4065
rect 12720 4045 12740 4065
rect 10470 3645 10490 3665
rect 10560 3645 10580 3665
rect 10650 3645 10670 3665
rect 10740 3645 10760 3665
rect 10830 3645 10850 3665
rect 10920 3645 10940 3665
rect 11010 3645 11030 3665
rect 11100 3645 11120 3665
rect 11190 3645 11210 3665
rect 11280 3645 11300 3665
rect 11370 3645 11390 3665
rect 11460 3645 11480 3665
rect 11550 3645 11570 3665
rect 11640 3645 11660 3665
rect 11730 3645 11750 3665
rect 11820 3645 11840 3665
rect 11910 3645 11930 3665
rect 12000 3645 12020 3665
rect 12090 3645 12110 3665
rect 12180 3645 12200 3665
rect 12270 3645 12290 3665
rect 12360 3645 12380 3665
rect 12450 3645 12470 3665
rect 12540 3645 12560 3665
rect 12630 3645 12650 3665
rect 12720 3645 12740 3665
rect 10470 3425 10490 3445
rect 10560 3425 10580 3445
rect 10650 3425 10670 3445
rect 10740 3425 10760 3445
rect 10830 3425 10850 3445
rect 10920 3425 10940 3445
rect 11010 3425 11030 3445
rect 11100 3425 11120 3445
rect 11190 3425 11210 3445
rect 11280 3425 11300 3445
rect 11370 3425 11390 3445
rect 11460 3425 11480 3445
rect 11550 3425 11570 3445
rect 11640 3425 11660 3445
rect 11730 3425 11750 3445
rect 11820 3425 11840 3445
rect 11910 3425 11930 3445
rect 12000 3425 12020 3445
rect 12090 3425 12110 3445
rect 12180 3425 12200 3445
rect 12270 3425 12290 3445
rect 12360 3425 12380 3445
rect 12450 3425 12470 3445
rect 12540 3425 12560 3445
rect 12630 3425 12650 3445
rect 12720 3425 12740 3445
<< nsubdiffcont >>
rect 10470 4345 10490 4365
rect 10560 4345 10580 4365
rect 10650 4345 10670 4365
rect 10740 4345 10760 4365
rect 10830 4345 10850 4365
rect 10920 4345 10940 4365
rect 11010 4345 11030 4365
rect 11100 4345 11120 4365
rect 11190 4345 11210 4365
rect 11280 4345 11300 4365
rect 11370 4345 11390 4365
rect 11460 4345 11480 4365
rect 11550 4345 11570 4365
rect 11640 4345 11660 4365
rect 11730 4345 11750 4365
rect 11820 4345 11840 4365
rect 11910 4345 11930 4365
rect 12000 4345 12020 4365
rect 12090 4345 12110 4365
rect 12180 4345 12200 4365
rect 12270 4345 12290 4365
rect 12360 4345 12380 4365
rect 12450 4345 12470 4365
rect 12540 4345 12560 4365
rect 12630 4345 12650 4365
rect 12720 4345 12740 4365
rect 10470 4125 10490 4145
rect 10560 4125 10580 4145
rect 10650 4125 10670 4145
rect 10740 4125 10760 4145
rect 10830 4125 10850 4145
rect 10920 4125 10940 4145
rect 11010 4125 11030 4145
rect 11100 4125 11120 4145
rect 11190 4125 11210 4145
rect 11280 4125 11300 4145
rect 11370 4125 11390 4145
rect 11460 4125 11480 4145
rect 11550 4125 11570 4145
rect 11640 4125 11660 4145
rect 11730 4125 11750 4145
rect 11820 4125 11840 4145
rect 11910 4125 11930 4145
rect 12000 4125 12020 4145
rect 12090 4125 12110 4145
rect 12180 4125 12200 4145
rect 12270 4125 12290 4145
rect 12360 4125 12380 4145
rect 12450 4125 12470 4145
rect 12540 4125 12560 4145
rect 12630 4125 12650 4145
rect 12720 4125 12740 4145
<< poly >>
rect 10455 4315 10505 4330
rect 10545 4315 10595 4330
rect 10635 4315 10685 4330
rect 10725 4315 10775 4330
rect 10815 4315 10865 4330
rect 10905 4315 10955 4330
rect 10995 4315 11045 4330
rect 11085 4315 11135 4330
rect 11175 4315 11225 4330
rect 11265 4315 11315 4330
rect 11355 4315 11405 4330
rect 11445 4315 11495 4330
rect 11535 4315 11585 4330
rect 11625 4315 11675 4330
rect 11715 4315 11765 4330
rect 11805 4315 11855 4330
rect 11895 4315 11945 4330
rect 11985 4315 12035 4330
rect 12075 4315 12125 4330
rect 12165 4315 12215 4330
rect 12255 4315 12305 4330
rect 12345 4315 12395 4330
rect 12435 4315 12485 4330
rect 12525 4315 12575 4330
rect 12615 4315 12665 4330
rect 12705 4315 12755 4330
rect 10455 4195 10505 4215
rect 10545 4195 10595 4215
rect 10455 4190 10595 4195
rect 10455 4170 10470 4190
rect 10490 4170 10560 4190
rect 10580 4170 10595 4190
rect 10455 4165 10595 4170
rect 10635 4195 10685 4215
rect 10725 4195 10775 4215
rect 10635 4190 10775 4195
rect 10635 4170 10650 4190
rect 10670 4170 10740 4190
rect 10760 4170 10775 4190
rect 10635 4165 10775 4170
rect 10815 4195 10865 4215
rect 10905 4195 10955 4215
rect 10815 4190 10955 4195
rect 10815 4170 10830 4190
rect 10850 4170 10920 4190
rect 10940 4170 10955 4190
rect 10815 4165 10955 4170
rect 10995 4195 11045 4215
rect 11085 4195 11135 4215
rect 10995 4190 11135 4195
rect 10995 4170 11010 4190
rect 11030 4170 11100 4190
rect 11120 4170 11135 4190
rect 10995 4165 11135 4170
rect 11175 4195 11225 4215
rect 11265 4195 11315 4215
rect 11175 4190 11315 4195
rect 11175 4170 11190 4190
rect 11210 4170 11280 4190
rect 11300 4170 11315 4190
rect 11175 4165 11315 4170
rect 11355 4195 11405 4215
rect 11445 4195 11495 4215
rect 11355 4190 11495 4195
rect 11355 4170 11370 4190
rect 11390 4170 11460 4190
rect 11480 4170 11495 4190
rect 11355 4165 11495 4170
rect 11535 4195 11585 4215
rect 11625 4195 11675 4215
rect 11535 4190 11675 4195
rect 11535 4170 11550 4190
rect 11570 4170 11640 4190
rect 11660 4170 11675 4190
rect 11535 4165 11675 4170
rect 11715 4195 11765 4215
rect 11805 4195 11855 4215
rect 11715 4190 11855 4195
rect 11715 4170 11730 4190
rect 11750 4170 11820 4190
rect 11840 4170 11855 4190
rect 11715 4165 11855 4170
rect 11895 4195 11945 4215
rect 11985 4195 12035 4215
rect 11895 4190 12035 4195
rect 11895 4170 11910 4190
rect 11930 4170 12000 4190
rect 12020 4170 12035 4190
rect 11895 4165 12035 4170
rect 12075 4195 12125 4215
rect 12165 4195 12215 4215
rect 12075 4190 12215 4195
rect 12075 4170 12090 4190
rect 12110 4170 12180 4190
rect 12200 4170 12215 4190
rect 12075 4165 12215 4170
rect 12255 4195 12305 4215
rect 12345 4195 12395 4215
rect 12255 4190 12395 4195
rect 12255 4170 12270 4190
rect 12290 4170 12360 4190
rect 12380 4170 12395 4190
rect 12255 4165 12395 4170
rect 12435 4195 12485 4215
rect 12525 4195 12575 4215
rect 12435 4190 12575 4195
rect 12435 4170 12450 4190
rect 12470 4170 12540 4190
rect 12560 4170 12575 4190
rect 12435 4165 12575 4170
rect 12615 4195 12665 4215
rect 12705 4195 12755 4215
rect 12615 4190 12755 4195
rect 12615 4170 12630 4190
rect 12650 4170 12720 4190
rect 12740 4170 12755 4190
rect 12615 4165 12755 4170
rect 10455 3620 10595 3625
rect 10455 3600 10470 3620
rect 10490 3600 10560 3620
rect 10580 3600 10595 3620
rect 10455 3595 10595 3600
rect 10455 3575 10505 3595
rect 10545 3575 10595 3595
rect 10635 3620 10775 3625
rect 10635 3600 10650 3620
rect 10670 3600 10740 3620
rect 10760 3600 10775 3620
rect 10635 3595 10775 3600
rect 10635 3575 10685 3595
rect 10725 3575 10775 3595
rect 10815 3620 10955 3625
rect 10815 3600 10830 3620
rect 10850 3600 10920 3620
rect 10940 3600 10955 3620
rect 10815 3595 10955 3600
rect 10815 3575 10865 3595
rect 10905 3575 10955 3595
rect 10995 3620 11135 3625
rect 10995 3600 11010 3620
rect 11030 3600 11100 3620
rect 11120 3600 11135 3620
rect 10995 3595 11135 3600
rect 10995 3575 11045 3595
rect 11085 3575 11135 3595
rect 11175 3620 11315 3625
rect 11175 3600 11190 3620
rect 11210 3600 11280 3620
rect 11300 3600 11315 3620
rect 11175 3595 11315 3600
rect 11175 3575 11225 3595
rect 11265 3575 11315 3595
rect 11355 3620 11495 3625
rect 11355 3600 11370 3620
rect 11390 3600 11460 3620
rect 11480 3600 11495 3620
rect 11355 3595 11495 3600
rect 11355 3575 11405 3595
rect 11445 3575 11495 3595
rect 11535 3620 11675 3625
rect 11535 3600 11550 3620
rect 11570 3600 11640 3620
rect 11660 3600 11675 3620
rect 11535 3595 11675 3600
rect 11535 3575 11585 3595
rect 11625 3575 11675 3595
rect 11715 3620 11855 3625
rect 11715 3600 11730 3620
rect 11750 3600 11820 3620
rect 11840 3600 11855 3620
rect 11715 3595 11855 3600
rect 11715 3575 11765 3595
rect 11805 3575 11855 3595
rect 11895 3620 12035 3625
rect 11895 3600 11910 3620
rect 11930 3600 12000 3620
rect 12020 3600 12035 3620
rect 11895 3595 12035 3600
rect 11895 3575 11945 3595
rect 11985 3575 12035 3595
rect 12075 3620 12215 3625
rect 12075 3600 12090 3620
rect 12110 3600 12180 3620
rect 12200 3600 12215 3620
rect 12075 3595 12215 3600
rect 12075 3575 12125 3595
rect 12165 3575 12215 3595
rect 12255 3620 12395 3625
rect 12255 3600 12270 3620
rect 12290 3600 12360 3620
rect 12380 3600 12395 3620
rect 12255 3595 12395 3600
rect 12255 3575 12305 3595
rect 12345 3575 12395 3595
rect 12435 3620 12575 3625
rect 12435 3600 12450 3620
rect 12470 3600 12540 3620
rect 12560 3600 12575 3620
rect 12435 3595 12575 3600
rect 12435 3575 12485 3595
rect 12525 3575 12575 3595
rect 12615 3620 12755 3625
rect 12615 3600 12630 3620
rect 12650 3600 12720 3620
rect 12740 3600 12755 3620
rect 12615 3595 12755 3600
rect 12615 3575 12665 3595
rect 12705 3575 12755 3595
rect 10455 3460 10505 3475
rect 10545 3460 10595 3475
rect 10635 3460 10685 3475
rect 10725 3460 10775 3475
rect 10815 3460 10865 3475
rect 10905 3460 10955 3475
rect 10995 3460 11045 3475
rect 11085 3460 11135 3475
rect 11175 3460 11225 3475
rect 11265 3460 11315 3475
rect 11355 3460 11405 3475
rect 11445 3460 11495 3475
rect 11535 3460 11585 3475
rect 11625 3460 11675 3475
rect 11715 3460 11765 3475
rect 11805 3460 11855 3475
rect 11895 3460 11945 3475
rect 11985 3460 12035 3475
rect 12075 3460 12125 3475
rect 12165 3460 12215 3475
rect 12255 3460 12305 3475
rect 12345 3460 12395 3475
rect 12435 3460 12485 3475
rect 12525 3460 12575 3475
rect 12615 3460 12665 3475
rect 12705 3460 12755 3475
<< polycont >>
rect 10470 4170 10490 4190
rect 10560 4170 10580 4190
rect 10650 4170 10670 4190
rect 10740 4170 10760 4190
rect 10830 4170 10850 4190
rect 10920 4170 10940 4190
rect 11010 4170 11030 4190
rect 11100 4170 11120 4190
rect 11190 4170 11210 4190
rect 11280 4170 11300 4190
rect 11370 4170 11390 4190
rect 11460 4170 11480 4190
rect 11550 4170 11570 4190
rect 11640 4170 11660 4190
rect 11730 4170 11750 4190
rect 11820 4170 11840 4190
rect 11910 4170 11930 4190
rect 12000 4170 12020 4190
rect 12090 4170 12110 4190
rect 12180 4170 12200 4190
rect 12270 4170 12290 4190
rect 12360 4170 12380 4190
rect 12450 4170 12470 4190
rect 12540 4170 12560 4190
rect 12630 4170 12650 4190
rect 12720 4170 12740 4190
rect 10470 3600 10490 3620
rect 10560 3600 10580 3620
rect 10650 3600 10670 3620
rect 10740 3600 10760 3620
rect 10830 3600 10850 3620
rect 10920 3600 10940 3620
rect 11010 3600 11030 3620
rect 11100 3600 11120 3620
rect 11190 3600 11210 3620
rect 11280 3600 11300 3620
rect 11370 3600 11390 3620
rect 11460 3600 11480 3620
rect 11550 3600 11570 3620
rect 11640 3600 11660 3620
rect 11730 3600 11750 3620
rect 11820 3600 11840 3620
rect 11910 3600 11930 3620
rect 12000 3600 12020 3620
rect 12090 3600 12110 3620
rect 12180 3600 12200 3620
rect 12270 3600 12290 3620
rect 12360 3600 12380 3620
rect 12450 3600 12470 3620
rect 12540 3600 12560 3620
rect 12630 3600 12650 3620
rect 12720 3600 12740 3620
<< locali >>
rect 10290 4065 10310 4375
rect 10365 4345 10425 4365
rect 10445 4345 10470 4365
rect 10490 4345 10560 4365
rect 10580 4345 10605 4365
rect 10625 4345 10650 4365
rect 10670 4345 10740 4365
rect 10760 4345 10785 4365
rect 10805 4345 10830 4365
rect 10850 4345 10920 4365
rect 10940 4345 10965 4365
rect 10985 4345 11010 4365
rect 11030 4345 11100 4365
rect 11120 4345 11145 4365
rect 11165 4345 11190 4365
rect 11210 4345 11280 4365
rect 11300 4345 11325 4365
rect 11345 4345 11370 4365
rect 11390 4345 11460 4365
rect 11480 4345 11505 4365
rect 11525 4345 11550 4365
rect 11570 4345 11640 4365
rect 11660 4345 11685 4365
rect 11705 4345 11730 4365
rect 11750 4345 11820 4365
rect 11840 4345 11865 4365
rect 11885 4345 11910 4365
rect 11930 4345 12000 4365
rect 12020 4345 12045 4365
rect 12065 4345 12090 4365
rect 12110 4345 12180 4365
rect 12200 4345 12225 4365
rect 12245 4345 12270 4365
rect 12290 4345 12360 4365
rect 12380 4345 12405 4365
rect 12425 4345 12450 4365
rect 12470 4345 12540 4365
rect 12560 4345 12585 4365
rect 12605 4345 12630 4365
rect 12650 4345 12720 4365
rect 12740 4345 12765 4365
rect 12785 4345 12794 4365
rect 10365 4145 10385 4345
rect 10425 4305 10445 4315
rect 10425 4215 10445 4225
rect 10515 4305 10535 4315
rect 10515 4190 10535 4225
rect 10605 4305 10625 4315
rect 10605 4215 10625 4225
rect 10695 4305 10715 4315
rect 10695 4215 10715 4225
rect 10785 4305 10805 4315
rect 10785 4215 10805 4225
rect 10875 4305 10895 4315
rect 10875 4215 10895 4225
rect 10965 4305 10985 4315
rect 10965 4215 10985 4225
rect 11055 4305 11075 4315
rect 11055 4215 11075 4225
rect 11145 4305 11165 4315
rect 11145 4215 11165 4225
rect 11235 4305 11255 4315
rect 11235 4215 11255 4225
rect 11325 4305 11345 4315
rect 11325 4215 11345 4225
rect 11415 4305 11435 4315
rect 11415 4215 11435 4225
rect 11505 4305 11525 4315
rect 11505 4215 11525 4225
rect 11595 4305 11615 4315
rect 11595 4215 11615 4225
rect 11685 4305 11705 4315
rect 11685 4215 11705 4225
rect 11775 4305 11795 4315
rect 11775 4215 11795 4225
rect 11865 4305 11885 4315
rect 11865 4215 11885 4225
rect 11955 4305 11975 4315
rect 11955 4215 11975 4225
rect 12045 4305 12065 4315
rect 12045 4215 12065 4225
rect 12135 4305 12155 4315
rect 12135 4215 12155 4225
rect 12225 4305 12245 4315
rect 12225 4215 12245 4225
rect 12315 4305 12335 4315
rect 12315 4215 12335 4225
rect 12405 4305 12425 4315
rect 12405 4215 12425 4225
rect 12495 4305 12515 4315
rect 12495 4215 12515 4225
rect 12585 4305 12605 4315
rect 12585 4215 12605 4225
rect 12675 4305 12695 4315
rect 12675 4215 12695 4225
rect 12765 4305 12785 4315
rect 12765 4215 12785 4225
rect 10460 4170 10470 4190
rect 10490 4170 10560 4190
rect 10580 4170 10599 4190
rect 10640 4170 10650 4190
rect 10670 4170 10740 4190
rect 10760 4170 10770 4190
rect 10820 4170 10830 4190
rect 10850 4170 10920 4190
rect 10940 4170 10950 4190
rect 11000 4170 11010 4190
rect 11030 4170 11100 4190
rect 11120 4170 11130 4190
rect 11180 4170 11190 4190
rect 11210 4170 11280 4190
rect 11300 4170 11310 4190
rect 11360 4170 11370 4190
rect 11390 4170 11460 4190
rect 11480 4170 11490 4190
rect 11540 4170 11550 4190
rect 11570 4170 11640 4190
rect 11660 4170 11670 4190
rect 11720 4170 11730 4190
rect 11750 4170 11820 4190
rect 11840 4170 11850 4190
rect 11900 4170 11910 4190
rect 11930 4170 12000 4190
rect 12020 4170 12030 4190
rect 12080 4170 12090 4190
rect 12110 4170 12180 4190
rect 12200 4170 12210 4190
rect 12260 4170 12270 4190
rect 12290 4170 12360 4190
rect 12380 4170 12390 4190
rect 12440 4170 12450 4190
rect 12470 4170 12540 4190
rect 12560 4170 12570 4190
rect 12620 4170 12630 4190
rect 12650 4170 12720 4190
rect 12740 4170 12750 4190
rect 10365 4125 10470 4145
rect 10490 4125 10560 4145
rect 10580 4125 10650 4145
rect 10670 4125 10740 4145
rect 10760 4125 10830 4145
rect 10850 4125 10920 4145
rect 10940 4125 11010 4145
rect 11030 4125 11100 4145
rect 11120 4125 11190 4145
rect 11210 4125 11280 4145
rect 11300 4125 11370 4145
rect 11390 4125 11460 4145
rect 11480 4125 11550 4145
rect 11570 4125 11640 4145
rect 11660 4125 11730 4145
rect 11750 4125 11820 4145
rect 11840 4125 11910 4145
rect 11930 4125 12000 4145
rect 12020 4125 12090 4145
rect 12110 4125 12180 4145
rect 12200 4125 12270 4145
rect 12290 4125 12360 4145
rect 12380 4125 12450 4145
rect 12470 4125 12540 4145
rect 12560 4125 12630 4145
rect 12650 4125 12720 4145
rect 12740 4125 12794 4145
rect 10415 4085 11370 4105
rect 11390 4085 11595 4105
rect 11615 4085 11685 4105
rect 11705 4085 11775 4105
rect 11795 4085 11910 4105
rect 11930 4085 12090 4105
rect 12110 4085 12630 4105
rect 12650 4085 12794 4105
rect 10290 4045 10470 4065
rect 10490 4045 10560 4065
rect 10580 4045 10650 4065
rect 10670 4045 10740 4065
rect 10760 4045 10830 4065
rect 10850 4045 10920 4065
rect 10940 4045 11010 4065
rect 11030 4045 11100 4065
rect 11120 4045 11190 4065
rect 11210 4045 11280 4065
rect 11300 4045 11370 4065
rect 11390 4045 11460 4065
rect 11480 4045 11550 4065
rect 11570 4045 11640 4065
rect 11660 4045 11730 4065
rect 11750 4045 11820 4065
rect 11840 4045 11910 4065
rect 11930 4045 12000 4065
rect 12020 4045 12090 4065
rect 12110 4045 12180 4065
rect 12200 4045 12270 4065
rect 12290 4045 12360 4065
rect 12380 4045 12450 4065
rect 12470 4045 12540 4065
rect 12560 4045 12630 4065
rect 12650 4045 12720 4065
rect 12740 4045 12794 4065
rect 10415 4005 11460 4025
rect 11480 4005 12000 4025
rect 12020 4005 12794 4025
rect 10415 3965 11640 3985
rect 11660 3965 11820 3985
rect 11840 3965 12794 3985
rect 10415 3925 10785 3945
rect 10805 3925 10965 3945
rect 10985 3925 11145 3945
rect 11165 3925 12225 3945
rect 12245 3925 12405 3945
rect 12425 3925 12585 3945
rect 12605 3925 12794 3945
rect 10415 3885 12270 3905
rect 12290 3885 12315 3905
rect 12335 3885 12360 3905
rect 12380 3885 12450 3905
rect 12470 3885 12495 3905
rect 12515 3885 12540 3905
rect 12560 3885 12794 3905
rect 10415 3845 10920 3865
rect 10940 3845 11100 3865
rect 11120 3845 11550 3865
rect 11570 3845 11730 3865
rect 11750 3845 12794 3865
rect 10415 3805 11505 3825
rect 11525 3805 11685 3825
rect 11705 3805 11865 3825
rect 11885 3805 12225 3825
rect 12245 3805 12405 3825
rect 12425 3805 12585 3825
rect 12605 3805 12794 3825
rect 10415 3765 10740 3785
rect 10760 3765 10875 3785
rect 10895 3765 10965 3785
rect 10985 3765 11055 3785
rect 11075 3765 11280 3785
rect 11300 3765 12180 3785
rect 12200 3765 12720 3785
rect 12740 3765 12794 3785
rect 10415 3725 10830 3745
rect 10850 3725 11010 3745
rect 11030 3725 12794 3745
rect 10415 3685 10650 3705
rect 10670 3685 11190 3705
rect 11210 3685 12794 3705
rect 10290 3645 10470 3665
rect 10490 3645 10560 3665
rect 10580 3645 10650 3665
rect 10670 3645 10740 3665
rect 10760 3645 10830 3665
rect 10850 3645 10920 3665
rect 10940 3645 11010 3665
rect 11030 3645 11100 3665
rect 11120 3645 11190 3665
rect 11210 3645 11280 3665
rect 11300 3645 11370 3665
rect 11390 3645 11460 3665
rect 11480 3645 11550 3665
rect 11570 3645 11640 3665
rect 11660 3645 11730 3665
rect 11750 3645 11820 3665
rect 11840 3645 11910 3665
rect 11930 3645 12000 3665
rect 12020 3645 12090 3665
rect 12110 3645 12180 3665
rect 12200 3645 12270 3665
rect 12290 3645 12360 3665
rect 12380 3645 12450 3665
rect 12470 3645 12540 3665
rect 12560 3645 12630 3665
rect 12650 3645 12720 3665
rect 12740 3645 12794 3665
rect 10290 3445 10310 3645
rect 10460 3600 10470 3620
rect 10490 3600 10560 3620
rect 10580 3600 10599 3620
rect 10640 3600 10650 3620
rect 10670 3600 10740 3620
rect 10760 3600 10770 3620
rect 10820 3600 10830 3620
rect 10850 3600 10920 3620
rect 10940 3600 10950 3620
rect 11000 3600 11010 3620
rect 11030 3600 11100 3620
rect 11120 3600 11130 3620
rect 11180 3600 11190 3620
rect 11210 3600 11280 3620
rect 11300 3600 11310 3620
rect 11360 3600 11370 3620
rect 11390 3600 11460 3620
rect 11480 3600 11490 3620
rect 11540 3600 11550 3620
rect 11570 3600 11640 3620
rect 11660 3600 11670 3620
rect 11720 3600 11730 3620
rect 11750 3600 11820 3620
rect 11840 3600 11850 3620
rect 11900 3600 11910 3620
rect 11930 3600 12000 3620
rect 12020 3600 12030 3620
rect 12080 3600 12090 3620
rect 12110 3600 12180 3620
rect 12200 3600 12210 3620
rect 12260 3600 12270 3620
rect 12290 3600 12360 3620
rect 12380 3600 12390 3620
rect 12440 3600 12450 3620
rect 12470 3600 12540 3620
rect 12560 3600 12570 3620
rect 12620 3600 12630 3620
rect 12650 3600 12720 3620
rect 12740 3600 12750 3620
rect 10425 3565 10445 3575
rect 10425 3475 10445 3485
rect 10515 3565 10535 3600
rect 10515 3475 10535 3485
rect 10605 3565 10625 3575
rect 10605 3475 10625 3485
rect 10695 3565 10715 3575
rect 10695 3475 10715 3485
rect 10785 3565 10805 3575
rect 10785 3475 10805 3485
rect 10875 3565 10895 3575
rect 10875 3475 10895 3485
rect 10965 3565 10985 3575
rect 10965 3475 10985 3485
rect 11055 3565 11075 3575
rect 11055 3475 11075 3485
rect 11145 3565 11165 3575
rect 11145 3475 11165 3485
rect 11235 3565 11255 3575
rect 11235 3475 11255 3485
rect 11325 3565 11345 3575
rect 11325 3475 11345 3485
rect 11415 3565 11435 3575
rect 11415 3475 11435 3485
rect 11505 3565 11525 3575
rect 11505 3475 11525 3485
rect 11595 3565 11615 3575
rect 11595 3475 11615 3485
rect 11685 3565 11705 3575
rect 11685 3475 11705 3485
rect 11775 3565 11795 3575
rect 11775 3475 11795 3485
rect 11865 3565 11885 3575
rect 11865 3475 11885 3485
rect 11955 3565 11975 3575
rect 11955 3475 11975 3485
rect 12045 3565 12065 3575
rect 12045 3475 12065 3485
rect 12135 3565 12155 3575
rect 12135 3475 12155 3485
rect 12225 3565 12245 3575
rect 12225 3475 12245 3485
rect 12315 3565 12335 3575
rect 12315 3475 12335 3485
rect 12405 3565 12425 3575
rect 12405 3475 12425 3485
rect 12495 3565 12515 3575
rect 12495 3475 12515 3485
rect 12585 3565 12605 3575
rect 12585 3475 12605 3485
rect 12675 3565 12695 3575
rect 12675 3475 12695 3485
rect 12765 3565 12785 3575
rect 12765 3475 12785 3485
rect 10280 3425 10290 3445
rect 10310 3425 10425 3445
rect 10445 3425 10470 3445
rect 10490 3425 10560 3445
rect 10580 3425 10605 3445
rect 10625 3425 10650 3445
rect 10670 3425 10740 3445
rect 10760 3425 10785 3445
rect 10805 3425 10830 3445
rect 10850 3425 10920 3445
rect 10940 3425 10965 3445
rect 10985 3425 11010 3445
rect 11030 3425 11100 3445
rect 11120 3425 11145 3445
rect 11165 3425 11190 3445
rect 11210 3425 11280 3445
rect 11300 3425 11325 3445
rect 11345 3425 11370 3445
rect 11390 3425 11460 3445
rect 11480 3425 11505 3445
rect 11525 3425 11550 3445
rect 11570 3425 11640 3445
rect 11660 3425 11685 3445
rect 11705 3425 11730 3445
rect 11750 3425 11820 3445
rect 11840 3425 11865 3445
rect 11885 3425 11910 3445
rect 11930 3425 12000 3445
rect 12020 3425 12045 3445
rect 12065 3425 12090 3445
rect 12110 3425 12180 3445
rect 12200 3425 12225 3445
rect 12245 3425 12270 3445
rect 12290 3425 12360 3445
rect 12380 3425 12405 3445
rect 12425 3425 12450 3445
rect 12470 3425 12540 3445
rect 12560 3425 12585 3445
rect 12605 3425 12630 3445
rect 12650 3425 12720 3445
rect 12740 3425 12765 3445
rect 12785 3425 12794 3445
<< viali >>
rect 10425 4345 10445 4365
rect 10605 4345 10625 4365
rect 10785 4345 10805 4365
rect 10965 4345 10985 4365
rect 11145 4345 11165 4365
rect 11325 4345 11345 4365
rect 11505 4345 11525 4365
rect 11685 4345 11705 4365
rect 11865 4345 11885 4365
rect 12045 4345 12065 4365
rect 12225 4345 12245 4365
rect 12405 4345 12425 4365
rect 12585 4345 12605 4365
rect 12765 4345 12785 4365
rect 10425 4225 10445 4305
rect 10605 4225 10625 4305
rect 10695 4225 10715 4305
rect 10785 4225 10805 4305
rect 10875 4225 10895 4305
rect 10965 4225 10985 4305
rect 11055 4225 11075 4305
rect 11145 4225 11165 4305
rect 11235 4225 11255 4305
rect 11325 4225 11345 4305
rect 11415 4225 11435 4305
rect 11505 4225 11525 4305
rect 11595 4225 11615 4305
rect 11685 4225 11705 4305
rect 11775 4225 11795 4305
rect 11865 4225 11885 4305
rect 11955 4225 11975 4305
rect 12045 4225 12065 4305
rect 12135 4225 12155 4305
rect 12225 4225 12245 4305
rect 12315 4225 12335 4305
rect 12405 4225 12425 4305
rect 12495 4225 12515 4305
rect 12585 4225 12605 4305
rect 12675 4225 12695 4305
rect 12765 4225 12785 4305
rect 10740 4170 10760 4190
rect 10920 4170 10940 4190
rect 11100 4170 11120 4190
rect 11280 4170 11300 4190
rect 11460 4170 11480 4190
rect 11640 4170 11660 4190
rect 11820 4170 11840 4190
rect 12000 4170 12020 4190
rect 12180 4170 12200 4190
rect 12360 4170 12380 4190
rect 12540 4170 12560 4190
rect 12720 4170 12740 4190
rect 11370 4085 11390 4105
rect 11595 4085 11615 4105
rect 11685 4085 11705 4105
rect 11775 4085 11795 4105
rect 11910 4085 11930 4105
rect 12090 4085 12110 4105
rect 12630 4085 12650 4105
rect 11460 4005 11480 4025
rect 12000 4005 12020 4025
rect 11640 3965 11660 3985
rect 11820 3965 11840 3985
rect 10785 3925 10805 3945
rect 10965 3925 10985 3945
rect 11145 3925 11165 3945
rect 12225 3925 12245 3945
rect 12405 3925 12425 3945
rect 12585 3925 12605 3945
rect 12270 3885 12290 3905
rect 12315 3885 12335 3905
rect 12360 3885 12380 3905
rect 12450 3885 12470 3905
rect 12495 3885 12515 3905
rect 12540 3885 12560 3905
rect 10920 3845 10940 3865
rect 11100 3845 11120 3865
rect 11550 3845 11570 3865
rect 11730 3845 11750 3865
rect 11505 3805 11525 3825
rect 11685 3805 11705 3825
rect 11865 3805 11885 3825
rect 12225 3805 12245 3825
rect 12405 3805 12425 3825
rect 12585 3805 12605 3825
rect 10740 3765 10760 3785
rect 10875 3765 10895 3785
rect 10965 3765 10985 3785
rect 11055 3765 11075 3785
rect 11280 3765 11300 3785
rect 12180 3765 12200 3785
rect 12720 3765 12740 3785
rect 10830 3725 10850 3745
rect 11010 3725 11030 3745
rect 10650 3685 10670 3705
rect 11190 3685 11210 3705
rect 10650 3600 10670 3620
rect 10830 3600 10850 3620
rect 11010 3600 11030 3620
rect 11190 3600 11210 3620
rect 11370 3600 11390 3620
rect 11550 3600 11570 3620
rect 11730 3600 11750 3620
rect 11910 3600 11930 3620
rect 12090 3600 12110 3620
rect 12270 3600 12290 3620
rect 12450 3600 12470 3620
rect 12630 3600 12650 3620
rect 10425 3485 10445 3565
rect 10605 3485 10625 3565
rect 10695 3485 10715 3565
rect 10785 3485 10805 3565
rect 10875 3485 10895 3565
rect 10965 3485 10985 3565
rect 11055 3485 11075 3565
rect 11145 3485 11165 3565
rect 11235 3485 11255 3565
rect 11325 3485 11345 3565
rect 11415 3485 11435 3565
rect 11505 3485 11525 3565
rect 11595 3485 11615 3565
rect 11685 3485 11705 3565
rect 11775 3485 11795 3565
rect 11865 3485 11885 3565
rect 11955 3485 11975 3565
rect 12045 3485 12065 3565
rect 12135 3485 12155 3565
rect 12225 3485 12245 3565
rect 12315 3485 12335 3565
rect 12405 3485 12425 3565
rect 12495 3485 12515 3565
rect 12585 3485 12605 3565
rect 12675 3485 12695 3565
rect 12765 3485 12785 3565
rect 10290 3425 10310 3445
rect 10425 3425 10445 3445
rect 10605 3425 10625 3445
rect 10785 3425 10805 3445
rect 10965 3425 10985 3445
rect 11145 3425 11165 3445
rect 11325 3425 11345 3445
rect 11505 3425 11525 3445
rect 11685 3425 11705 3445
rect 11865 3425 11885 3445
rect 12045 3425 12065 3445
rect 12225 3425 12245 3445
rect 12405 3425 12425 3445
rect 12585 3425 12605 3445
rect 12765 3425 12785 3445
<< metal1 >>
rect 10280 3450 10320 4375
rect 10415 4370 10455 4375
rect 10415 4340 10420 4370
rect 10450 4340 10455 4370
rect 10415 4335 10455 4340
rect 10425 4315 10445 4335
rect 10515 4315 10535 4375
rect 10596 4370 10635 4375
rect 10596 4340 10600 4370
rect 10630 4340 10635 4370
rect 10596 4335 10635 4340
rect 10775 4370 10815 4375
rect 10775 4340 10780 4370
rect 10810 4340 10815 4370
rect 10775 4335 10815 4340
rect 10955 4370 10995 4375
rect 10955 4340 10960 4370
rect 10990 4340 10995 4370
rect 10955 4335 10995 4340
rect 11135 4370 11175 4375
rect 11135 4340 11140 4370
rect 11170 4340 11175 4370
rect 11135 4335 11175 4340
rect 11315 4370 11355 4375
rect 11315 4340 11320 4370
rect 11350 4340 11355 4370
rect 11315 4335 11355 4340
rect 11495 4370 11535 4375
rect 11495 4340 11500 4370
rect 11530 4340 11535 4370
rect 11495 4335 11535 4340
rect 11675 4370 11715 4375
rect 11675 4340 11680 4370
rect 11710 4340 11715 4370
rect 11675 4335 11715 4340
rect 11855 4370 11895 4375
rect 11855 4340 11860 4370
rect 11890 4340 11895 4370
rect 11855 4335 11895 4340
rect 12035 4370 12075 4375
rect 12035 4340 12040 4370
rect 12070 4340 12075 4370
rect 12035 4335 12075 4340
rect 12215 4370 12255 4375
rect 12215 4340 12220 4370
rect 12250 4340 12255 4370
rect 12215 4335 12255 4340
rect 12395 4370 12435 4375
rect 12395 4340 12400 4370
rect 12430 4340 12435 4370
rect 12395 4335 12435 4340
rect 12575 4370 12615 4375
rect 12575 4340 12580 4370
rect 12610 4340 12615 4370
rect 12575 4335 12615 4340
rect 12755 4370 12794 4375
rect 12755 4340 12760 4370
rect 12790 4340 12794 4370
rect 12755 4335 12794 4340
rect 10605 4315 10625 4335
rect 11325 4315 11345 4335
rect 12045 4315 12065 4335
rect 12765 4315 12785 4335
rect 10420 4305 10450 4315
rect 10420 4225 10425 4305
rect 10445 4225 10450 4305
rect 10420 4215 10450 4225
rect 10510 4215 10540 4315
rect 10600 4305 10630 4315
rect 10600 4225 10605 4305
rect 10625 4225 10630 4305
rect 10600 4215 10630 4225
rect 10690 4305 10720 4315
rect 10690 4225 10695 4305
rect 10715 4225 10720 4305
rect 10690 4215 10720 4225
rect 10780 4305 10810 4315
rect 10780 4225 10785 4305
rect 10805 4225 10810 4305
rect 10780 4215 10810 4225
rect 10870 4305 10900 4315
rect 10870 4225 10875 4305
rect 10895 4225 10900 4305
rect 10870 4215 10900 4225
rect 10960 4305 10990 4315
rect 10960 4225 10965 4305
rect 10985 4225 10990 4305
rect 10960 4215 10990 4225
rect 11050 4305 11080 4315
rect 11050 4225 11055 4305
rect 11075 4225 11080 4305
rect 11050 4215 11080 4225
rect 11140 4305 11170 4315
rect 11140 4225 11145 4305
rect 11165 4225 11170 4305
rect 11140 4215 11170 4225
rect 11230 4305 11260 4315
rect 11230 4225 11235 4305
rect 11255 4225 11260 4305
rect 11230 4215 11260 4225
rect 11320 4305 11350 4315
rect 11320 4225 11325 4305
rect 11345 4225 11350 4305
rect 11320 4215 11350 4225
rect 11410 4305 11440 4315
rect 11410 4225 11415 4305
rect 11435 4225 11440 4305
rect 11410 4215 11440 4225
rect 11500 4305 11530 4315
rect 11500 4225 11505 4305
rect 11525 4225 11530 4305
rect 11500 4215 11530 4225
rect 11590 4305 11620 4315
rect 11590 4225 11595 4305
rect 11615 4225 11620 4305
rect 11590 4215 11620 4225
rect 11680 4305 11710 4315
rect 11680 4225 11685 4305
rect 11705 4225 11710 4305
rect 11680 4215 11710 4225
rect 11770 4305 11800 4315
rect 11770 4225 11775 4305
rect 11795 4225 11800 4305
rect 11770 4215 11800 4225
rect 11860 4305 11890 4315
rect 11860 4225 11865 4305
rect 11885 4225 11890 4305
rect 11860 4215 11890 4225
rect 11950 4305 11980 4315
rect 11950 4225 11955 4305
rect 11975 4225 11980 4305
rect 11950 4215 11980 4225
rect 12040 4305 12070 4315
rect 12040 4225 12045 4305
rect 12065 4225 12070 4305
rect 12040 4215 12070 4225
rect 12130 4305 12160 4315
rect 12130 4225 12135 4305
rect 12155 4225 12160 4305
rect 12130 4215 12160 4225
rect 12220 4305 12250 4315
rect 12220 4225 12225 4305
rect 12245 4225 12250 4305
rect 12220 4215 12250 4225
rect 12310 4305 12340 4315
rect 12310 4225 12315 4305
rect 12335 4225 12340 4305
rect 12310 4215 12340 4225
rect 12400 4305 12430 4315
rect 12400 4225 12405 4305
rect 12425 4225 12430 4305
rect 12400 4215 12430 4225
rect 12490 4305 12520 4315
rect 12490 4225 12495 4305
rect 12515 4225 12520 4305
rect 12490 4215 12520 4225
rect 12580 4305 12610 4315
rect 12580 4225 12585 4305
rect 12605 4225 12610 4305
rect 12580 4215 12610 4225
rect 12670 4305 12700 4315
rect 12670 4225 12675 4305
rect 12695 4225 12700 4305
rect 12670 4215 12700 4225
rect 12760 4305 12790 4315
rect 12760 4225 12765 4305
rect 12785 4225 12790 4305
rect 12760 4215 12790 4225
rect 10515 3575 10535 4215
rect 10740 4195 10760 4200
rect 10735 4190 10765 4195
rect 10735 4170 10740 4190
rect 10760 4170 10765 4190
rect 10735 4165 10765 4170
rect 10740 3790 10760 4165
rect 10785 3950 10805 4215
rect 10780 3945 10810 3950
rect 10780 3925 10785 3945
rect 10805 3925 10810 3945
rect 10780 3920 10810 3925
rect 10785 3915 10805 3920
rect 10875 3790 10895 4215
rect 10920 4195 10940 4200
rect 10915 4190 10945 4195
rect 10915 4170 10920 4190
rect 10940 4170 10945 4190
rect 10915 4165 10945 4170
rect 10920 3870 10940 4165
rect 10965 3950 10985 4215
rect 10960 3945 10990 3950
rect 10960 3925 10965 3945
rect 10985 3925 10990 3945
rect 10960 3920 10990 3925
rect 10965 3915 10985 3920
rect 10915 3865 10945 3870
rect 10915 3845 10920 3865
rect 10940 3845 10945 3865
rect 10915 3840 10945 3845
rect 10920 3835 10940 3840
rect 10965 3790 10985 3795
rect 11055 3790 11075 4215
rect 11100 4195 11120 4200
rect 11095 4190 11125 4195
rect 11095 4170 11100 4190
rect 11120 4170 11125 4190
rect 11095 4165 11125 4170
rect 11100 3870 11120 4165
rect 11145 3950 11165 4215
rect 11280 4195 11300 4200
rect 11460 4195 11480 4200
rect 11640 4195 11660 4200
rect 11275 4190 11305 4195
rect 11275 4170 11280 4190
rect 11300 4170 11305 4190
rect 11275 4165 11305 4170
rect 11455 4190 11485 4195
rect 11455 4170 11460 4190
rect 11480 4170 11485 4190
rect 11455 4165 11485 4170
rect 11635 4190 11665 4195
rect 11635 4170 11640 4190
rect 11660 4170 11665 4190
rect 11635 4165 11665 4170
rect 11140 3945 11170 3950
rect 11140 3925 11145 3945
rect 11165 3925 11170 3945
rect 11140 3920 11170 3925
rect 11145 3915 11165 3920
rect 11095 3865 11125 3870
rect 11095 3845 11100 3865
rect 11120 3845 11125 3865
rect 11095 3840 11125 3845
rect 11100 3835 11120 3840
rect 11280 3790 11300 4165
rect 11370 4110 11390 4115
rect 11365 4105 11395 4110
rect 11365 4085 11370 4105
rect 11390 4085 11395 4105
rect 11365 4080 11395 4085
rect 10735 3785 10765 3790
rect 10735 3765 10740 3785
rect 10760 3765 10765 3785
rect 10735 3760 10765 3765
rect 10870 3785 10900 3790
rect 10870 3765 10875 3785
rect 10895 3765 10900 3785
rect 10870 3760 10900 3765
rect 10960 3785 10990 3790
rect 10960 3765 10965 3785
rect 10985 3765 10990 3785
rect 10960 3760 10990 3765
rect 11050 3785 11080 3790
rect 11050 3765 11055 3785
rect 11075 3765 11080 3785
rect 11050 3760 11080 3765
rect 11275 3785 11305 3790
rect 11275 3765 11280 3785
rect 11300 3765 11305 3785
rect 11275 3760 11305 3765
rect 10740 3755 10760 3760
rect 10875 3755 10895 3760
rect 10830 3750 10850 3755
rect 10825 3745 10855 3750
rect 10825 3725 10830 3745
rect 10850 3725 10855 3745
rect 10825 3720 10855 3725
rect 10650 3710 10670 3715
rect 10645 3705 10675 3710
rect 10645 3685 10650 3705
rect 10670 3685 10675 3705
rect 10645 3680 10675 3685
rect 10650 3625 10670 3680
rect 10830 3625 10850 3720
rect 10645 3620 10675 3625
rect 10645 3600 10650 3620
rect 10670 3600 10675 3620
rect 10645 3595 10675 3600
rect 10825 3620 10855 3625
rect 10825 3600 10830 3620
rect 10850 3600 10855 3620
rect 10825 3595 10855 3600
rect 10650 3590 10670 3595
rect 10830 3590 10850 3595
rect 10605 3575 10625 3580
rect 10965 3575 10985 3760
rect 11055 3755 11075 3760
rect 11280 3755 11300 3760
rect 11010 3750 11030 3755
rect 11005 3745 11035 3750
rect 11005 3725 11010 3745
rect 11030 3725 11035 3745
rect 11005 3720 11035 3725
rect 11010 3625 11030 3720
rect 11190 3710 11210 3715
rect 11185 3705 11215 3710
rect 11185 3685 11190 3705
rect 11210 3685 11215 3705
rect 11185 3680 11215 3685
rect 11190 3625 11210 3680
rect 11370 3625 11390 4080
rect 11460 4030 11480 4165
rect 11595 4110 11615 4115
rect 11590 4105 11620 4110
rect 11590 4085 11595 4105
rect 11615 4085 11620 4105
rect 11590 4080 11620 4085
rect 11455 4025 11485 4030
rect 11455 4005 11460 4025
rect 11480 4005 11485 4025
rect 11455 4000 11485 4005
rect 11460 3995 11480 4000
rect 11550 3870 11570 3875
rect 11545 3865 11575 3870
rect 11545 3845 11550 3865
rect 11570 3845 11575 3865
rect 11545 3840 11575 3845
rect 11505 3830 11525 3835
rect 11500 3825 11530 3830
rect 11500 3805 11505 3825
rect 11525 3805 11530 3825
rect 11500 3800 11530 3805
rect 11005 3620 11035 3625
rect 11005 3600 11010 3620
rect 11030 3600 11035 3620
rect 11005 3595 11035 3600
rect 11185 3620 11215 3625
rect 11185 3600 11190 3620
rect 11210 3600 11215 3620
rect 11185 3595 11215 3600
rect 11365 3620 11395 3625
rect 11365 3600 11370 3620
rect 11390 3600 11395 3620
rect 11365 3595 11395 3600
rect 11010 3590 11030 3595
rect 11190 3590 11210 3595
rect 11370 3590 11390 3595
rect 11505 3575 11525 3800
rect 11550 3625 11570 3840
rect 11545 3620 11575 3625
rect 11545 3600 11550 3620
rect 11570 3600 11575 3620
rect 11545 3595 11575 3600
rect 11550 3590 11570 3595
rect 11595 3575 11615 4080
rect 11640 3990 11660 4165
rect 11685 4110 11705 4215
rect 11865 4210 11885 4215
rect 11820 4195 11840 4200
rect 12000 4195 12020 4200
rect 12180 4195 12200 4200
rect 11815 4190 11845 4195
rect 11815 4170 11820 4190
rect 11840 4170 11845 4190
rect 11815 4165 11845 4170
rect 11995 4190 12025 4195
rect 11995 4170 12000 4190
rect 12020 4170 12025 4190
rect 11995 4165 12025 4170
rect 12175 4190 12205 4195
rect 12175 4170 12180 4190
rect 12200 4170 12205 4190
rect 12175 4165 12205 4170
rect 11775 4110 11795 4115
rect 11680 4105 11710 4110
rect 11680 4085 11685 4105
rect 11705 4085 11710 4105
rect 11680 4080 11710 4085
rect 11770 4105 11800 4110
rect 11770 4085 11775 4105
rect 11795 4085 11800 4105
rect 11770 4080 11800 4085
rect 11685 4075 11705 4080
rect 11635 3985 11665 3990
rect 11635 3965 11640 3985
rect 11660 3965 11665 3985
rect 11635 3960 11665 3965
rect 11640 3955 11660 3960
rect 11730 3870 11750 3875
rect 11725 3865 11755 3870
rect 11725 3845 11730 3865
rect 11750 3845 11755 3865
rect 11725 3840 11755 3845
rect 11685 3830 11705 3835
rect 11680 3825 11710 3830
rect 11680 3805 11685 3825
rect 11705 3805 11710 3825
rect 11680 3800 11710 3805
rect 11685 3575 11705 3800
rect 11730 3625 11750 3840
rect 11725 3620 11755 3625
rect 11725 3600 11730 3620
rect 11750 3600 11755 3620
rect 11725 3595 11755 3600
rect 11730 3590 11750 3595
rect 11775 3575 11795 4080
rect 11820 3990 11840 4165
rect 11910 4110 11930 4115
rect 11905 4105 11935 4110
rect 11905 4085 11910 4105
rect 11930 4085 11935 4105
rect 11905 4080 11935 4085
rect 11815 3985 11845 3990
rect 11815 3965 11820 3985
rect 11840 3965 11845 3985
rect 11815 3960 11845 3965
rect 11820 3955 11840 3960
rect 11865 3830 11885 3835
rect 11860 3825 11890 3830
rect 11860 3805 11865 3825
rect 11885 3805 11890 3825
rect 11860 3800 11890 3805
rect 11865 3575 11885 3800
rect 11910 3625 11930 4080
rect 12000 4030 12020 4165
rect 12090 4110 12110 4115
rect 12085 4105 12115 4110
rect 12085 4085 12090 4105
rect 12110 4085 12115 4105
rect 12085 4080 12115 4085
rect 11995 4025 12025 4030
rect 11995 4005 12000 4025
rect 12020 4005 12025 4025
rect 11995 4000 12025 4005
rect 12000 3995 12020 4000
rect 12090 3625 12110 4080
rect 12180 3790 12200 4165
rect 12225 3950 12245 4215
rect 12220 3945 12250 3950
rect 12220 3925 12225 3945
rect 12245 3925 12250 3945
rect 12220 3920 12250 3925
rect 12225 3915 12245 3920
rect 12270 3910 12290 3915
rect 12315 3910 12335 4215
rect 12360 4195 12380 4200
rect 12355 4190 12385 4195
rect 12355 4170 12360 4190
rect 12380 4170 12385 4190
rect 12355 4165 12385 4170
rect 12360 3910 12380 4165
rect 12405 3950 12425 4215
rect 12400 3945 12430 3950
rect 12400 3925 12405 3945
rect 12425 3925 12430 3945
rect 12400 3920 12430 3925
rect 12405 3915 12425 3920
rect 12450 3910 12470 3915
rect 12495 3910 12515 4215
rect 12540 4195 12560 4200
rect 12535 4190 12565 4195
rect 12535 4170 12540 4190
rect 12560 4170 12565 4190
rect 12535 4165 12565 4170
rect 12540 3910 12560 4165
rect 12585 3950 12605 4215
rect 12720 4195 12740 4200
rect 12715 4190 12745 4195
rect 12715 4170 12720 4190
rect 12740 4170 12745 4190
rect 12715 4165 12745 4170
rect 12630 4110 12650 4115
rect 12625 4105 12655 4110
rect 12625 4085 12630 4105
rect 12650 4085 12655 4105
rect 12625 4080 12655 4085
rect 12580 3945 12610 3950
rect 12580 3925 12585 3945
rect 12605 3925 12610 3945
rect 12580 3920 12610 3925
rect 12585 3915 12605 3920
rect 12265 3905 12295 3910
rect 12265 3885 12270 3905
rect 12290 3885 12295 3905
rect 12265 3880 12295 3885
rect 12310 3905 12340 3910
rect 12310 3885 12315 3905
rect 12335 3885 12340 3905
rect 12310 3880 12340 3885
rect 12355 3905 12385 3910
rect 12355 3885 12360 3905
rect 12380 3885 12385 3905
rect 12355 3880 12385 3885
rect 12445 3905 12475 3910
rect 12445 3885 12450 3905
rect 12470 3885 12475 3905
rect 12445 3880 12475 3885
rect 12490 3905 12520 3910
rect 12490 3885 12495 3905
rect 12515 3885 12520 3905
rect 12490 3880 12520 3885
rect 12535 3905 12565 3910
rect 12535 3885 12540 3905
rect 12560 3885 12565 3905
rect 12535 3880 12565 3885
rect 12225 3830 12245 3835
rect 12220 3825 12250 3830
rect 12220 3805 12225 3825
rect 12245 3805 12250 3825
rect 12220 3800 12250 3805
rect 12175 3785 12205 3790
rect 12175 3765 12180 3785
rect 12200 3765 12205 3785
rect 12175 3760 12205 3765
rect 12180 3755 12200 3760
rect 11905 3620 11935 3625
rect 11905 3600 11910 3620
rect 11930 3600 11935 3620
rect 11905 3595 11935 3600
rect 12085 3620 12115 3625
rect 12085 3600 12090 3620
rect 12110 3600 12115 3620
rect 12085 3595 12115 3600
rect 11910 3590 11930 3595
rect 12090 3590 12110 3595
rect 12225 3575 12245 3800
rect 12270 3625 12290 3880
rect 12265 3620 12295 3625
rect 12265 3600 12270 3620
rect 12290 3600 12295 3620
rect 12265 3595 12295 3600
rect 12270 3590 12290 3595
rect 12315 3575 12335 3880
rect 12360 3875 12380 3880
rect 12405 3830 12425 3835
rect 12400 3825 12430 3830
rect 12400 3805 12405 3825
rect 12425 3805 12430 3825
rect 12400 3800 12430 3805
rect 12405 3575 12425 3800
rect 12450 3625 12470 3880
rect 12445 3620 12475 3625
rect 12445 3600 12450 3620
rect 12470 3600 12475 3620
rect 12445 3595 12475 3600
rect 12450 3590 12470 3595
rect 12495 3575 12515 3880
rect 12540 3875 12560 3880
rect 12585 3830 12605 3835
rect 12580 3825 12610 3830
rect 12580 3805 12585 3825
rect 12605 3805 12610 3825
rect 12580 3800 12610 3805
rect 12585 3575 12605 3800
rect 12630 3625 12650 4080
rect 12720 3790 12740 4165
rect 12715 3785 12745 3790
rect 12715 3765 12720 3785
rect 12740 3765 12745 3785
rect 12715 3760 12745 3765
rect 12720 3755 12740 3760
rect 12625 3620 12655 3625
rect 12625 3600 12630 3620
rect 12650 3600 12655 3620
rect 12625 3595 12655 3600
rect 12630 3590 12650 3595
rect 10420 3565 10450 3575
rect 10420 3485 10425 3565
rect 10445 3485 10450 3565
rect 10420 3475 10450 3485
rect 10510 3475 10540 3575
rect 10600 3565 10630 3575
rect 10600 3485 10605 3565
rect 10625 3485 10630 3565
rect 10600 3475 10630 3485
rect 10690 3565 10720 3575
rect 10690 3485 10695 3565
rect 10715 3485 10720 3565
rect 10690 3475 10720 3485
rect 10780 3565 10810 3575
rect 10780 3485 10785 3565
rect 10805 3485 10810 3565
rect 10780 3475 10810 3485
rect 10870 3565 10900 3575
rect 10870 3485 10875 3565
rect 10895 3485 10900 3565
rect 10870 3475 10900 3485
rect 10960 3565 10990 3575
rect 10960 3485 10965 3565
rect 10985 3485 10990 3565
rect 10960 3475 10990 3485
rect 11050 3565 11080 3575
rect 11050 3485 11055 3565
rect 11075 3485 11080 3565
rect 11050 3475 11080 3485
rect 11140 3565 11170 3575
rect 11140 3485 11145 3565
rect 11165 3485 11170 3565
rect 11140 3475 11170 3485
rect 11230 3565 11260 3575
rect 11230 3485 11235 3565
rect 11255 3485 11260 3565
rect 11230 3475 11260 3485
rect 11320 3565 11350 3575
rect 11320 3485 11325 3565
rect 11345 3485 11350 3565
rect 11320 3475 11350 3485
rect 11410 3565 11440 3575
rect 11410 3485 11415 3565
rect 11435 3485 11440 3565
rect 11410 3475 11440 3485
rect 11500 3565 11530 3575
rect 11500 3485 11505 3565
rect 11525 3485 11530 3565
rect 11500 3475 11530 3485
rect 11590 3565 11620 3575
rect 11590 3485 11595 3565
rect 11615 3485 11620 3565
rect 11590 3475 11620 3485
rect 11680 3565 11710 3575
rect 11680 3485 11685 3565
rect 11705 3485 11710 3565
rect 11680 3475 11710 3485
rect 11770 3565 11800 3575
rect 11770 3485 11775 3565
rect 11795 3485 11800 3565
rect 11770 3475 11800 3485
rect 11860 3565 11890 3575
rect 11860 3485 11865 3565
rect 11885 3485 11890 3565
rect 11860 3475 11890 3485
rect 11950 3565 11980 3575
rect 11950 3485 11955 3565
rect 11975 3485 11980 3565
rect 11950 3475 11980 3485
rect 12040 3565 12070 3575
rect 12040 3485 12045 3565
rect 12065 3485 12070 3565
rect 12040 3475 12070 3485
rect 12130 3565 12160 3575
rect 12130 3485 12135 3565
rect 12155 3485 12160 3565
rect 12130 3475 12160 3485
rect 12220 3565 12250 3575
rect 12220 3485 12225 3565
rect 12245 3485 12250 3565
rect 12220 3475 12250 3485
rect 12310 3565 12340 3575
rect 12310 3485 12315 3565
rect 12335 3485 12340 3565
rect 12310 3475 12340 3485
rect 12400 3565 12430 3575
rect 12400 3485 12405 3565
rect 12425 3485 12430 3565
rect 12400 3475 12430 3485
rect 12490 3565 12520 3575
rect 12490 3485 12495 3565
rect 12515 3485 12520 3565
rect 12490 3475 12520 3485
rect 12580 3565 12610 3575
rect 12580 3485 12585 3565
rect 12605 3485 12610 3565
rect 12580 3475 12610 3485
rect 12670 3565 12700 3575
rect 12670 3485 12675 3565
rect 12695 3485 12700 3565
rect 12670 3475 12700 3485
rect 12760 3565 12790 3575
rect 12760 3485 12765 3565
rect 12785 3485 12790 3565
rect 12760 3475 12790 3485
rect 10425 3455 10445 3475
rect 10605 3455 10625 3475
rect 11325 3455 11345 3475
rect 12045 3455 12065 3475
rect 12765 3455 12785 3475
rect 10280 3420 10285 3450
rect 10315 3420 10320 3450
rect 10280 3415 10320 3420
rect 10415 3450 10455 3455
rect 10415 3420 10420 3450
rect 10450 3420 10455 3450
rect 10415 3415 10455 3420
rect 10596 3450 10635 3455
rect 10596 3420 10600 3450
rect 10630 3420 10635 3450
rect 10596 3415 10635 3420
rect 10775 3450 10815 3455
rect 10775 3420 10780 3450
rect 10810 3420 10815 3450
rect 10775 3415 10815 3420
rect 10955 3450 10995 3455
rect 10955 3420 10960 3450
rect 10990 3420 10995 3450
rect 10955 3415 10995 3420
rect 11135 3450 11175 3455
rect 11135 3420 11140 3450
rect 11170 3420 11175 3450
rect 11135 3415 11175 3420
rect 11315 3450 11355 3455
rect 11315 3420 11320 3450
rect 11350 3420 11355 3450
rect 11315 3415 11355 3420
rect 11495 3450 11535 3455
rect 11495 3420 11500 3450
rect 11530 3420 11535 3450
rect 11495 3415 11535 3420
rect 11675 3450 11715 3455
rect 11675 3420 11680 3450
rect 11710 3420 11715 3450
rect 11675 3415 11715 3420
rect 11855 3450 11895 3455
rect 11855 3420 11860 3450
rect 11890 3420 11895 3450
rect 11855 3415 11895 3420
rect 12035 3450 12075 3455
rect 12035 3420 12040 3450
rect 12070 3420 12075 3450
rect 12035 3415 12075 3420
rect 12215 3450 12255 3455
rect 12215 3420 12220 3450
rect 12250 3420 12255 3450
rect 12215 3415 12255 3420
rect 12395 3450 12435 3455
rect 12395 3420 12400 3450
rect 12430 3420 12435 3450
rect 12395 3415 12435 3420
rect 12575 3450 12615 3455
rect 12575 3420 12580 3450
rect 12610 3420 12615 3450
rect 12575 3415 12615 3420
rect 12755 3450 12794 3455
rect 12755 3420 12760 3450
rect 12790 3420 12794 3450
rect 12755 3415 12794 3420
<< via1 >>
rect 10420 4365 10450 4370
rect 10420 4345 10425 4365
rect 10425 4345 10445 4365
rect 10445 4345 10450 4365
rect 10420 4340 10450 4345
rect 10600 4365 10630 4370
rect 10600 4345 10605 4365
rect 10605 4345 10625 4365
rect 10625 4345 10630 4365
rect 10600 4340 10630 4345
rect 10780 4365 10810 4370
rect 10780 4345 10785 4365
rect 10785 4345 10805 4365
rect 10805 4345 10810 4365
rect 10780 4340 10810 4345
rect 10960 4365 10990 4370
rect 10960 4345 10965 4365
rect 10965 4345 10985 4365
rect 10985 4345 10990 4365
rect 10960 4340 10990 4345
rect 11140 4365 11170 4370
rect 11140 4345 11145 4365
rect 11145 4345 11165 4365
rect 11165 4345 11170 4365
rect 11140 4340 11170 4345
rect 11320 4365 11350 4370
rect 11320 4345 11325 4365
rect 11325 4345 11345 4365
rect 11345 4345 11350 4365
rect 11320 4340 11350 4345
rect 11500 4365 11530 4370
rect 11500 4345 11505 4365
rect 11505 4345 11525 4365
rect 11525 4345 11530 4365
rect 11500 4340 11530 4345
rect 11680 4365 11710 4370
rect 11680 4345 11685 4365
rect 11685 4345 11705 4365
rect 11705 4345 11710 4365
rect 11680 4340 11710 4345
rect 11860 4365 11890 4370
rect 11860 4345 11865 4365
rect 11865 4345 11885 4365
rect 11885 4345 11890 4365
rect 11860 4340 11890 4345
rect 12040 4365 12070 4370
rect 12040 4345 12045 4365
rect 12045 4345 12065 4365
rect 12065 4345 12070 4365
rect 12040 4340 12070 4345
rect 12220 4365 12250 4370
rect 12220 4345 12225 4365
rect 12225 4345 12245 4365
rect 12245 4345 12250 4365
rect 12220 4340 12250 4345
rect 12400 4365 12430 4370
rect 12400 4345 12405 4365
rect 12405 4345 12425 4365
rect 12425 4345 12430 4365
rect 12400 4340 12430 4345
rect 12580 4365 12610 4370
rect 12580 4345 12585 4365
rect 12585 4345 12605 4365
rect 12605 4345 12610 4365
rect 12580 4340 12610 4345
rect 12760 4365 12790 4370
rect 12760 4345 12765 4365
rect 12765 4345 12785 4365
rect 12785 4345 12790 4365
rect 12760 4340 12790 4345
rect 10285 3445 10315 3450
rect 10285 3425 10290 3445
rect 10290 3425 10310 3445
rect 10310 3425 10315 3445
rect 10285 3420 10315 3425
rect 10420 3445 10450 3450
rect 10420 3425 10425 3445
rect 10425 3425 10445 3445
rect 10445 3425 10450 3445
rect 10420 3420 10450 3425
rect 10600 3445 10630 3450
rect 10600 3425 10605 3445
rect 10605 3425 10625 3445
rect 10625 3425 10630 3445
rect 10600 3420 10630 3425
rect 10780 3445 10810 3450
rect 10780 3425 10785 3445
rect 10785 3425 10805 3445
rect 10805 3425 10810 3445
rect 10780 3420 10810 3425
rect 10960 3445 10990 3450
rect 10960 3425 10965 3445
rect 10965 3425 10985 3445
rect 10985 3425 10990 3445
rect 10960 3420 10990 3425
rect 11140 3445 11170 3450
rect 11140 3425 11145 3445
rect 11145 3425 11165 3445
rect 11165 3425 11170 3445
rect 11140 3420 11170 3425
rect 11320 3445 11350 3450
rect 11320 3425 11325 3445
rect 11325 3425 11345 3445
rect 11345 3425 11350 3445
rect 11320 3420 11350 3425
rect 11500 3445 11530 3450
rect 11500 3425 11505 3445
rect 11505 3425 11525 3445
rect 11525 3425 11530 3445
rect 11500 3420 11530 3425
rect 11680 3445 11710 3450
rect 11680 3425 11685 3445
rect 11685 3425 11705 3445
rect 11705 3425 11710 3445
rect 11680 3420 11710 3425
rect 11860 3445 11890 3450
rect 11860 3425 11865 3445
rect 11865 3425 11885 3445
rect 11885 3425 11890 3445
rect 11860 3420 11890 3425
rect 12040 3445 12070 3450
rect 12040 3425 12045 3445
rect 12045 3425 12065 3445
rect 12065 3425 12070 3445
rect 12040 3420 12070 3425
rect 12220 3445 12250 3450
rect 12220 3425 12225 3445
rect 12225 3425 12245 3445
rect 12245 3425 12250 3445
rect 12220 3420 12250 3425
rect 12400 3445 12430 3450
rect 12400 3425 12405 3445
rect 12405 3425 12425 3445
rect 12425 3425 12430 3445
rect 12400 3420 12430 3425
rect 12580 3445 12610 3450
rect 12580 3425 12585 3445
rect 12585 3425 12605 3445
rect 12605 3425 12610 3445
rect 12580 3420 12610 3425
rect 12760 3445 12790 3450
rect 12760 3425 12765 3445
rect 12765 3425 12785 3445
rect 12785 3425 12790 3445
rect 12760 3420 12790 3425
<< metal2 >>
rect 10415 4370 12794 4375
rect 10415 4340 10420 4370
rect 10450 4340 10600 4370
rect 10630 4340 10780 4370
rect 10810 4340 10960 4370
rect 10990 4340 11140 4370
rect 11170 4340 11320 4370
rect 11350 4340 11500 4370
rect 11530 4340 11680 4370
rect 11710 4340 11860 4370
rect 11890 4340 12040 4370
rect 12070 4340 12220 4370
rect 12250 4340 12400 4370
rect 12430 4340 12580 4370
rect 12610 4340 12760 4370
rect 12790 4340 12794 4370
rect 10415 4335 12794 4340
rect 10280 3450 12794 3455
rect 10280 3420 10285 3450
rect 10315 3420 10420 3450
rect 10450 3420 10600 3450
rect 10630 3420 10780 3450
rect 10810 3420 10960 3450
rect 10990 3420 11140 3450
rect 11170 3420 11320 3450
rect 11350 3420 11500 3450
rect 11530 3420 11680 3450
rect 11710 3420 11860 3450
rect 11890 3420 12040 3450
rect 12070 3420 12220 3450
rect 12250 3420 12400 3450
rect 12430 3420 12580 3450
rect 12610 3420 12760 3450
rect 12790 3420 12794 3450
rect 10280 3415 12794 3420
<< labels >>
rlabel locali 10425 3815 10425 3815 1 xn
rlabel locali 10425 3935 10425 3935 1 xp
rlabel locali 10425 4095 10425 4095 1 n3
rlabel locali 10425 3775 10425 3775 1 p3
rlabel locali 10425 3895 10425 3895 1 out
port 8 n
rlabel locali 10425 3735 10425 3735 1 n2
port 5 n
rlabel locali 10425 3695 10425 3695 1 n1
port 6 n
rlabel locali 10425 4015 10425 4015 1 p1
port 3 n
rlabel locali 10425 3975 10425 3975 1 p2
port 4 n
rlabel locali 10425 3855 10425 3855 1 in
port 7 n
rlabel metal2 10420 4355 10420 4355 1 VDDA
port 1 n
rlabel metal2 10420 3435 10420 3435 1 VSSA
port 2 n
<< end >>
