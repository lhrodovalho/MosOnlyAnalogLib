magic
tech sky130A
timestamp 1624076896
<< nwell >>
rect 9105 4375 20800 4385
rect 9105 4105 20805 4375
<< mvnmos >>
rect 9215 3475 9265 3575
rect 9305 3475 9355 3575
rect 9395 3475 9445 3575
rect 9485 3475 9535 3575
rect 9575 3475 9625 3575
rect 9665 3475 9715 3575
rect 9755 3475 9805 3575
rect 9845 3475 9895 3575
rect 9935 3475 9985 3575
rect 10025 3475 10075 3575
rect 10115 3475 10165 3575
rect 10205 3475 10255 3575
rect 10295 3475 10345 3575
rect 10385 3475 10435 3575
rect 10475 3475 10525 3575
rect 10565 3475 10615 3575
rect 10655 3475 10705 3575
rect 10745 3475 10795 3575
rect 10835 3475 10885 3575
rect 10925 3475 10975 3575
rect 11015 3475 11065 3575
rect 11105 3475 11155 3575
rect 11195 3475 11245 3575
rect 11285 3475 11335 3575
rect 11375 3475 11425 3575
rect 11465 3475 11515 3575
rect 11555 3475 11605 3575
rect 11645 3475 11695 3575
rect 11735 3475 11785 3575
rect 11825 3475 11875 3575
rect 11915 3475 11965 3575
rect 12005 3475 12055 3575
rect 12095 3475 12145 3575
rect 12185 3475 12235 3575
rect 12275 3475 12325 3575
rect 12365 3475 12415 3575
rect 12455 3475 12505 3575
rect 12545 3475 12595 3575
rect 12635 3475 12685 3575
rect 12725 3475 12775 3575
rect 12815 3475 12865 3575
rect 12905 3475 12955 3575
rect 12995 3475 13045 3575
rect 13085 3475 13135 3575
rect 13175 3475 13225 3575
rect 13265 3475 13315 3575
rect 13355 3475 13405 3575
rect 13445 3475 13495 3575
rect 13535 3475 13585 3575
rect 13625 3475 13675 3575
rect 13715 3475 13765 3575
rect 13805 3475 13855 3575
rect 13895 3475 13945 3575
rect 13985 3475 14035 3575
rect 14075 3475 14125 3575
rect 14165 3475 14215 3575
rect 14255 3475 14305 3575
rect 14345 3475 14395 3575
rect 14435 3475 14485 3575
rect 14525 3475 14575 3575
rect 14615 3475 14665 3575
rect 14705 3475 14755 3575
rect 14795 3475 14845 3575
rect 14885 3475 14935 3575
rect 14975 3475 15025 3575
rect 15065 3475 15115 3575
rect 15155 3475 15205 3575
rect 15245 3475 15295 3575
rect 15335 3475 15385 3575
rect 15425 3475 15475 3575
rect 15515 3475 15565 3575
rect 15605 3475 15655 3575
rect 15695 3475 15745 3575
rect 15785 3475 15835 3575
rect 15875 3475 15925 3575
rect 15965 3475 16015 3575
rect 16055 3475 16105 3575
rect 16145 3475 16195 3575
rect 16235 3475 16285 3575
rect 16325 3475 16375 3575
rect 16415 3475 16465 3575
rect 16505 3475 16555 3575
rect 16595 3475 16645 3575
rect 16685 3475 16735 3575
rect 16775 3475 16825 3575
rect 16865 3475 16915 3575
rect 16955 3475 17005 3575
rect 17045 3475 17095 3575
rect 17135 3475 17185 3575
rect 17225 3475 17275 3575
rect 17315 3475 17365 3575
rect 17405 3475 17455 3575
rect 17495 3475 17545 3575
rect 17585 3475 17635 3575
rect 17675 3475 17725 3575
rect 17765 3475 17815 3575
rect 17855 3475 17905 3575
rect 17945 3475 17995 3575
rect 18035 3475 18085 3575
rect 18125 3475 18175 3575
rect 18215 3475 18265 3575
rect 18305 3475 18355 3575
rect 18395 3475 18445 3575
rect 18485 3475 18535 3575
rect 18575 3475 18625 3575
rect 18665 3475 18715 3575
rect 18755 3475 18805 3575
rect 18845 3475 18895 3575
rect 18935 3475 18985 3575
rect 19025 3475 19075 3575
rect 19115 3475 19165 3575
rect 19205 3475 19255 3575
rect 19295 3475 19345 3575
rect 19385 3475 19435 3575
rect 19475 3475 19525 3575
rect 19565 3475 19615 3575
rect 19655 3475 19705 3575
rect 19745 3475 19795 3575
rect 19835 3475 19885 3575
rect 19925 3475 19975 3575
rect 20015 3475 20065 3575
rect 20105 3475 20155 3575
rect 20195 3475 20245 3575
rect 20285 3475 20335 3575
rect 20375 3475 20425 3575
rect 20465 3475 20515 3575
rect 20555 3475 20605 3575
rect 20645 3475 20695 3575
<< mvpmos >>
rect 9215 4215 9265 4315
rect 9305 4215 9355 4315
rect 9395 4215 9445 4315
rect 9485 4215 9535 4315
rect 9575 4215 9625 4315
rect 9665 4215 9715 4315
rect 9755 4215 9805 4315
rect 9845 4215 9895 4315
rect 9935 4215 9985 4315
rect 10025 4215 10075 4315
rect 10115 4215 10165 4315
rect 10205 4215 10255 4315
rect 10295 4215 10345 4315
rect 10385 4215 10435 4315
rect 10475 4215 10525 4315
rect 10565 4215 10615 4315
rect 10655 4215 10705 4315
rect 10745 4215 10795 4315
rect 10835 4215 10885 4315
rect 10925 4215 10975 4315
rect 11015 4215 11065 4315
rect 11105 4215 11155 4315
rect 11195 4215 11245 4315
rect 11285 4215 11335 4315
rect 11375 4215 11425 4315
rect 11465 4215 11515 4315
rect 11555 4215 11605 4315
rect 11645 4215 11695 4315
rect 11735 4215 11785 4315
rect 11825 4215 11875 4315
rect 11915 4215 11965 4315
rect 12005 4215 12055 4315
rect 12095 4215 12145 4315
rect 12185 4215 12235 4315
rect 12275 4215 12325 4315
rect 12365 4215 12415 4315
rect 12455 4215 12505 4315
rect 12545 4215 12595 4315
rect 12635 4215 12685 4315
rect 12725 4215 12775 4315
rect 12815 4215 12865 4315
rect 12905 4215 12955 4315
rect 12995 4215 13045 4315
rect 13085 4215 13135 4315
rect 13175 4215 13225 4315
rect 13265 4215 13315 4315
rect 13355 4215 13405 4315
rect 13445 4215 13495 4315
rect 13535 4215 13585 4315
rect 13625 4215 13675 4315
rect 13715 4215 13765 4315
rect 13805 4215 13855 4315
rect 13895 4215 13945 4315
rect 13985 4215 14035 4315
rect 14075 4215 14125 4315
rect 14165 4215 14215 4315
rect 14255 4215 14305 4315
rect 14345 4215 14395 4315
rect 14435 4215 14485 4315
rect 14525 4215 14575 4315
rect 14615 4215 14665 4315
rect 14705 4215 14755 4315
rect 14795 4215 14845 4315
rect 14885 4215 14935 4315
rect 14975 4215 15025 4315
rect 15065 4215 15115 4315
rect 15155 4215 15205 4315
rect 15245 4215 15295 4315
rect 15335 4215 15385 4315
rect 15425 4215 15475 4315
rect 15515 4215 15565 4315
rect 15605 4215 15655 4315
rect 15695 4215 15745 4315
rect 15785 4215 15835 4315
rect 15875 4215 15925 4315
rect 15965 4215 16015 4315
rect 16055 4215 16105 4315
rect 16145 4215 16195 4315
rect 16235 4215 16285 4315
rect 16325 4215 16375 4315
rect 16415 4215 16465 4315
rect 16505 4215 16555 4315
rect 16595 4215 16645 4315
rect 16685 4215 16735 4315
rect 16775 4215 16825 4315
rect 16865 4215 16915 4315
rect 16955 4215 17005 4315
rect 17045 4215 17095 4315
rect 17135 4215 17185 4315
rect 17225 4215 17275 4315
rect 17315 4215 17365 4315
rect 17405 4215 17455 4315
rect 17495 4215 17545 4315
rect 17585 4215 17635 4315
rect 17675 4215 17725 4315
rect 17765 4215 17815 4315
rect 17855 4215 17905 4315
rect 17945 4215 17995 4315
rect 18035 4215 18085 4315
rect 18125 4215 18175 4315
rect 18215 4215 18265 4315
rect 18305 4215 18355 4315
rect 18395 4215 18445 4315
rect 18485 4215 18535 4315
rect 18575 4215 18625 4315
rect 18665 4215 18715 4315
rect 18755 4215 18805 4315
rect 18845 4215 18895 4315
rect 18935 4215 18985 4315
rect 19025 4215 19075 4315
rect 19115 4215 19165 4315
rect 19205 4215 19255 4315
rect 19295 4215 19345 4315
rect 19385 4215 19435 4315
rect 19475 4215 19525 4315
rect 19565 4215 19615 4315
rect 19655 4215 19705 4315
rect 19745 4215 19795 4315
rect 19835 4215 19885 4315
rect 19925 4215 19975 4315
rect 20015 4215 20065 4315
rect 20105 4215 20155 4315
rect 20195 4215 20245 4315
rect 20285 4215 20335 4315
rect 20375 4215 20425 4315
rect 20465 4215 20515 4315
rect 20555 4215 20605 4315
rect 20645 4215 20695 4315
<< mvndiff >>
rect 9175 3565 9215 3575
rect 9175 3485 9185 3565
rect 9205 3485 9215 3565
rect 9175 3475 9215 3485
rect 9265 3565 9305 3575
rect 9265 3485 9275 3565
rect 9295 3485 9305 3565
rect 9265 3475 9305 3485
rect 9355 3565 9395 3575
rect 9355 3485 9365 3565
rect 9385 3485 9395 3565
rect 9355 3475 9395 3485
rect 9445 3565 9485 3575
rect 9445 3485 9455 3565
rect 9475 3485 9485 3565
rect 9445 3475 9485 3485
rect 9535 3565 9575 3575
rect 9535 3485 9545 3565
rect 9565 3485 9575 3565
rect 9535 3475 9575 3485
rect 9625 3565 9665 3575
rect 9625 3485 9635 3565
rect 9655 3485 9665 3565
rect 9625 3475 9665 3485
rect 9715 3565 9755 3575
rect 9715 3485 9725 3565
rect 9745 3485 9755 3565
rect 9715 3475 9755 3485
rect 9805 3565 9845 3575
rect 9805 3485 9815 3565
rect 9835 3485 9845 3565
rect 9805 3475 9845 3485
rect 9895 3565 9935 3575
rect 9895 3485 9905 3565
rect 9925 3485 9935 3565
rect 9895 3475 9935 3485
rect 9985 3565 10025 3575
rect 9985 3485 9995 3565
rect 10015 3485 10025 3565
rect 9985 3475 10025 3485
rect 10075 3565 10115 3575
rect 10075 3485 10085 3565
rect 10105 3485 10115 3565
rect 10075 3475 10115 3485
rect 10165 3565 10205 3575
rect 10165 3485 10175 3565
rect 10195 3485 10205 3565
rect 10165 3475 10205 3485
rect 10255 3565 10295 3575
rect 10255 3485 10265 3565
rect 10285 3485 10295 3565
rect 10255 3475 10295 3485
rect 10345 3565 10385 3575
rect 10345 3485 10355 3565
rect 10375 3485 10385 3565
rect 10345 3475 10385 3485
rect 10435 3565 10475 3575
rect 10435 3485 10445 3565
rect 10465 3485 10475 3565
rect 10435 3475 10475 3485
rect 10525 3565 10565 3575
rect 10525 3485 10535 3565
rect 10555 3485 10565 3565
rect 10525 3475 10565 3485
rect 10615 3565 10655 3575
rect 10615 3485 10625 3565
rect 10645 3485 10655 3565
rect 10615 3475 10655 3485
rect 10705 3565 10745 3575
rect 10705 3485 10715 3565
rect 10735 3485 10745 3565
rect 10705 3475 10745 3485
rect 10795 3565 10835 3575
rect 10795 3485 10805 3565
rect 10825 3485 10835 3565
rect 10795 3475 10835 3485
rect 10885 3565 10925 3575
rect 10885 3485 10895 3565
rect 10915 3485 10925 3565
rect 10885 3475 10925 3485
rect 10975 3565 11015 3575
rect 10975 3485 10985 3565
rect 11005 3485 11015 3565
rect 10975 3475 11015 3485
rect 11065 3565 11105 3575
rect 11065 3485 11075 3565
rect 11095 3485 11105 3565
rect 11065 3475 11105 3485
rect 11155 3565 11195 3575
rect 11155 3485 11165 3565
rect 11185 3485 11195 3565
rect 11155 3475 11195 3485
rect 11245 3565 11285 3575
rect 11245 3485 11255 3565
rect 11275 3485 11285 3565
rect 11245 3475 11285 3485
rect 11335 3565 11375 3575
rect 11335 3485 11345 3565
rect 11365 3485 11375 3565
rect 11335 3475 11375 3485
rect 11425 3565 11465 3575
rect 11425 3485 11435 3565
rect 11455 3485 11465 3565
rect 11425 3475 11465 3485
rect 11515 3565 11555 3575
rect 11515 3485 11525 3565
rect 11545 3485 11555 3565
rect 11515 3475 11555 3485
rect 11605 3565 11645 3575
rect 11605 3485 11615 3565
rect 11635 3485 11645 3565
rect 11605 3475 11645 3485
rect 11695 3565 11735 3575
rect 11695 3485 11705 3565
rect 11725 3485 11735 3565
rect 11695 3475 11735 3485
rect 11785 3565 11825 3575
rect 11785 3485 11795 3565
rect 11815 3485 11825 3565
rect 11785 3475 11825 3485
rect 11875 3565 11915 3575
rect 11875 3485 11885 3565
rect 11905 3485 11915 3565
rect 11875 3475 11915 3485
rect 11965 3565 12005 3575
rect 11965 3485 11975 3565
rect 11995 3485 12005 3565
rect 11965 3475 12005 3485
rect 12055 3565 12095 3575
rect 12055 3485 12065 3565
rect 12085 3485 12095 3565
rect 12055 3475 12095 3485
rect 12145 3565 12185 3575
rect 12145 3485 12155 3565
rect 12175 3485 12185 3565
rect 12145 3475 12185 3485
rect 12235 3565 12275 3575
rect 12235 3485 12245 3565
rect 12265 3485 12275 3565
rect 12235 3475 12275 3485
rect 12325 3565 12365 3575
rect 12325 3485 12335 3565
rect 12355 3485 12365 3565
rect 12325 3475 12365 3485
rect 12415 3565 12455 3575
rect 12415 3485 12425 3565
rect 12445 3485 12455 3565
rect 12415 3475 12455 3485
rect 12505 3565 12545 3575
rect 12505 3485 12515 3565
rect 12535 3485 12545 3565
rect 12505 3475 12545 3485
rect 12595 3565 12635 3575
rect 12595 3485 12605 3565
rect 12625 3485 12635 3565
rect 12595 3475 12635 3485
rect 12685 3565 12725 3575
rect 12685 3485 12695 3565
rect 12715 3485 12725 3565
rect 12685 3475 12725 3485
rect 12775 3565 12815 3575
rect 12775 3485 12785 3565
rect 12805 3485 12815 3565
rect 12775 3475 12815 3485
rect 12865 3565 12905 3575
rect 12865 3485 12875 3565
rect 12895 3485 12905 3565
rect 12865 3475 12905 3485
rect 12955 3565 12995 3575
rect 12955 3485 12965 3565
rect 12985 3485 12995 3565
rect 12955 3475 12995 3485
rect 13045 3565 13085 3575
rect 13045 3485 13055 3565
rect 13075 3485 13085 3565
rect 13045 3475 13085 3485
rect 13135 3565 13175 3575
rect 13135 3485 13145 3565
rect 13165 3485 13175 3565
rect 13135 3475 13175 3485
rect 13225 3565 13265 3575
rect 13225 3485 13235 3565
rect 13255 3485 13265 3565
rect 13225 3475 13265 3485
rect 13315 3565 13355 3575
rect 13315 3485 13325 3565
rect 13345 3485 13355 3565
rect 13315 3475 13355 3485
rect 13405 3565 13445 3575
rect 13405 3485 13415 3565
rect 13435 3485 13445 3565
rect 13405 3475 13445 3485
rect 13495 3565 13535 3575
rect 13495 3485 13505 3565
rect 13525 3485 13535 3565
rect 13495 3475 13535 3485
rect 13585 3565 13625 3575
rect 13585 3485 13595 3565
rect 13615 3485 13625 3565
rect 13585 3475 13625 3485
rect 13675 3565 13715 3575
rect 13675 3485 13685 3565
rect 13705 3485 13715 3565
rect 13675 3475 13715 3485
rect 13765 3565 13805 3575
rect 13765 3485 13775 3565
rect 13795 3485 13805 3565
rect 13765 3475 13805 3485
rect 13855 3565 13895 3575
rect 13855 3485 13865 3565
rect 13885 3485 13895 3565
rect 13855 3475 13895 3485
rect 13945 3565 13985 3575
rect 13945 3485 13955 3565
rect 13975 3485 13985 3565
rect 13945 3475 13985 3485
rect 14035 3565 14075 3575
rect 14035 3485 14045 3565
rect 14065 3485 14075 3565
rect 14035 3475 14075 3485
rect 14125 3565 14165 3575
rect 14125 3485 14135 3565
rect 14155 3485 14165 3565
rect 14125 3475 14165 3485
rect 14215 3565 14255 3575
rect 14215 3485 14225 3565
rect 14245 3485 14255 3565
rect 14215 3475 14255 3485
rect 14305 3565 14345 3575
rect 14305 3485 14315 3565
rect 14335 3485 14345 3565
rect 14305 3475 14345 3485
rect 14395 3565 14435 3575
rect 14395 3485 14405 3565
rect 14425 3485 14435 3565
rect 14395 3475 14435 3485
rect 14485 3565 14525 3575
rect 14485 3485 14495 3565
rect 14515 3485 14525 3565
rect 14485 3475 14525 3485
rect 14575 3565 14615 3575
rect 14575 3485 14585 3565
rect 14605 3485 14615 3565
rect 14575 3475 14615 3485
rect 14665 3565 14705 3575
rect 14665 3485 14675 3565
rect 14695 3485 14705 3565
rect 14665 3475 14705 3485
rect 14755 3565 14795 3575
rect 14755 3485 14765 3565
rect 14785 3485 14795 3565
rect 14755 3475 14795 3485
rect 14845 3565 14885 3575
rect 14845 3485 14855 3565
rect 14875 3485 14885 3565
rect 14845 3475 14885 3485
rect 14935 3565 14975 3575
rect 14935 3485 14945 3565
rect 14965 3485 14975 3565
rect 14935 3475 14975 3485
rect 15025 3565 15065 3575
rect 15025 3485 15035 3565
rect 15055 3485 15065 3565
rect 15025 3475 15065 3485
rect 15115 3565 15155 3575
rect 15115 3485 15125 3565
rect 15145 3485 15155 3565
rect 15115 3475 15155 3485
rect 15205 3565 15245 3575
rect 15205 3485 15215 3565
rect 15235 3485 15245 3565
rect 15205 3475 15245 3485
rect 15295 3565 15335 3575
rect 15295 3485 15305 3565
rect 15325 3485 15335 3565
rect 15295 3475 15335 3485
rect 15385 3565 15425 3575
rect 15385 3485 15395 3565
rect 15415 3485 15425 3565
rect 15385 3475 15425 3485
rect 15475 3565 15515 3575
rect 15475 3485 15485 3565
rect 15505 3485 15515 3565
rect 15475 3475 15515 3485
rect 15565 3565 15605 3575
rect 15565 3485 15575 3565
rect 15595 3485 15605 3565
rect 15565 3475 15605 3485
rect 15655 3565 15695 3575
rect 15655 3485 15665 3565
rect 15685 3485 15695 3565
rect 15655 3475 15695 3485
rect 15745 3565 15785 3575
rect 15745 3485 15755 3565
rect 15775 3485 15785 3565
rect 15745 3475 15785 3485
rect 15835 3565 15875 3575
rect 15835 3485 15845 3565
rect 15865 3485 15875 3565
rect 15835 3475 15875 3485
rect 15925 3565 15965 3575
rect 15925 3485 15935 3565
rect 15955 3485 15965 3565
rect 15925 3475 15965 3485
rect 16015 3565 16055 3575
rect 16015 3485 16025 3565
rect 16045 3485 16055 3565
rect 16015 3475 16055 3485
rect 16105 3565 16145 3575
rect 16105 3485 16115 3565
rect 16135 3485 16145 3565
rect 16105 3475 16145 3485
rect 16195 3565 16235 3575
rect 16195 3485 16205 3565
rect 16225 3485 16235 3565
rect 16195 3475 16235 3485
rect 16285 3565 16325 3575
rect 16285 3485 16295 3565
rect 16315 3485 16325 3565
rect 16285 3475 16325 3485
rect 16375 3565 16415 3575
rect 16375 3485 16385 3565
rect 16405 3485 16415 3565
rect 16375 3475 16415 3485
rect 16465 3565 16505 3575
rect 16465 3485 16475 3565
rect 16495 3485 16505 3565
rect 16465 3475 16505 3485
rect 16555 3565 16595 3575
rect 16555 3485 16565 3565
rect 16585 3485 16595 3565
rect 16555 3475 16595 3485
rect 16645 3565 16685 3575
rect 16645 3485 16655 3565
rect 16675 3485 16685 3565
rect 16645 3475 16685 3485
rect 16735 3565 16775 3575
rect 16735 3485 16745 3565
rect 16765 3485 16775 3565
rect 16735 3475 16775 3485
rect 16825 3565 16865 3575
rect 16825 3485 16835 3565
rect 16855 3485 16865 3565
rect 16825 3475 16865 3485
rect 16915 3565 16955 3575
rect 16915 3485 16925 3565
rect 16945 3485 16955 3565
rect 16915 3475 16955 3485
rect 17005 3565 17045 3575
rect 17005 3485 17015 3565
rect 17035 3485 17045 3565
rect 17005 3475 17045 3485
rect 17095 3565 17135 3575
rect 17095 3485 17105 3565
rect 17125 3485 17135 3565
rect 17095 3475 17135 3485
rect 17185 3565 17225 3575
rect 17185 3485 17195 3565
rect 17215 3485 17225 3565
rect 17185 3475 17225 3485
rect 17275 3565 17315 3575
rect 17275 3485 17285 3565
rect 17305 3485 17315 3565
rect 17275 3475 17315 3485
rect 17365 3565 17405 3575
rect 17365 3485 17375 3565
rect 17395 3485 17405 3565
rect 17365 3475 17405 3485
rect 17455 3565 17495 3575
rect 17455 3485 17465 3565
rect 17485 3485 17495 3565
rect 17455 3475 17495 3485
rect 17545 3565 17585 3575
rect 17545 3485 17555 3565
rect 17575 3485 17585 3565
rect 17545 3475 17585 3485
rect 17635 3565 17675 3575
rect 17635 3485 17645 3565
rect 17665 3485 17675 3565
rect 17635 3475 17675 3485
rect 17725 3565 17765 3575
rect 17725 3485 17735 3565
rect 17755 3485 17765 3565
rect 17725 3475 17765 3485
rect 17815 3565 17855 3575
rect 17815 3485 17825 3565
rect 17845 3485 17855 3565
rect 17815 3475 17855 3485
rect 17905 3565 17945 3575
rect 17905 3485 17915 3565
rect 17935 3485 17945 3565
rect 17905 3475 17945 3485
rect 17995 3565 18035 3575
rect 17995 3485 18005 3565
rect 18025 3485 18035 3565
rect 17995 3475 18035 3485
rect 18085 3565 18125 3575
rect 18085 3485 18095 3565
rect 18115 3485 18125 3565
rect 18085 3475 18125 3485
rect 18175 3565 18215 3575
rect 18175 3485 18185 3565
rect 18205 3485 18215 3565
rect 18175 3475 18215 3485
rect 18265 3565 18305 3575
rect 18265 3485 18275 3565
rect 18295 3485 18305 3565
rect 18265 3475 18305 3485
rect 18355 3565 18395 3575
rect 18355 3485 18365 3565
rect 18385 3485 18395 3565
rect 18355 3475 18395 3485
rect 18445 3565 18485 3575
rect 18445 3485 18455 3565
rect 18475 3485 18485 3565
rect 18445 3475 18485 3485
rect 18535 3565 18575 3575
rect 18535 3485 18545 3565
rect 18565 3485 18575 3565
rect 18535 3475 18575 3485
rect 18625 3565 18665 3575
rect 18625 3485 18635 3565
rect 18655 3485 18665 3565
rect 18625 3475 18665 3485
rect 18715 3565 18755 3575
rect 18715 3485 18725 3565
rect 18745 3485 18755 3565
rect 18715 3475 18755 3485
rect 18805 3565 18845 3575
rect 18805 3485 18815 3565
rect 18835 3485 18845 3565
rect 18805 3475 18845 3485
rect 18895 3565 18935 3575
rect 18895 3485 18905 3565
rect 18925 3485 18935 3565
rect 18895 3475 18935 3485
rect 18985 3565 19025 3575
rect 18985 3485 18995 3565
rect 19015 3485 19025 3565
rect 18985 3475 19025 3485
rect 19075 3565 19115 3575
rect 19075 3485 19085 3565
rect 19105 3485 19115 3565
rect 19075 3475 19115 3485
rect 19165 3565 19205 3575
rect 19165 3485 19175 3565
rect 19195 3485 19205 3565
rect 19165 3475 19205 3485
rect 19255 3565 19295 3575
rect 19255 3485 19265 3565
rect 19285 3485 19295 3565
rect 19255 3475 19295 3485
rect 19345 3565 19385 3575
rect 19345 3485 19355 3565
rect 19375 3485 19385 3565
rect 19345 3475 19385 3485
rect 19435 3565 19475 3575
rect 19435 3485 19445 3565
rect 19465 3485 19475 3565
rect 19435 3475 19475 3485
rect 19525 3565 19565 3575
rect 19525 3485 19535 3565
rect 19555 3485 19565 3565
rect 19525 3475 19565 3485
rect 19615 3565 19655 3575
rect 19615 3485 19625 3565
rect 19645 3485 19655 3565
rect 19615 3475 19655 3485
rect 19705 3565 19745 3575
rect 19705 3485 19715 3565
rect 19735 3485 19745 3565
rect 19705 3475 19745 3485
rect 19795 3565 19835 3575
rect 19795 3485 19805 3565
rect 19825 3485 19835 3565
rect 19795 3475 19835 3485
rect 19885 3565 19925 3575
rect 19885 3485 19895 3565
rect 19915 3485 19925 3565
rect 19885 3475 19925 3485
rect 19975 3565 20015 3575
rect 19975 3485 19985 3565
rect 20005 3485 20015 3565
rect 19975 3475 20015 3485
rect 20065 3565 20105 3575
rect 20065 3485 20075 3565
rect 20095 3485 20105 3565
rect 20065 3475 20105 3485
rect 20155 3565 20195 3575
rect 20155 3485 20165 3565
rect 20185 3485 20195 3565
rect 20155 3475 20195 3485
rect 20245 3565 20285 3575
rect 20245 3485 20255 3565
rect 20275 3485 20285 3565
rect 20245 3475 20285 3485
rect 20335 3565 20375 3575
rect 20335 3485 20345 3565
rect 20365 3485 20375 3565
rect 20335 3475 20375 3485
rect 20425 3565 20465 3575
rect 20425 3485 20435 3565
rect 20455 3485 20465 3565
rect 20425 3475 20465 3485
rect 20515 3565 20555 3575
rect 20515 3485 20525 3565
rect 20545 3485 20555 3565
rect 20515 3475 20555 3485
rect 20605 3565 20645 3575
rect 20605 3485 20615 3565
rect 20635 3485 20645 3565
rect 20605 3475 20645 3485
rect 20695 3565 20735 3575
rect 20695 3485 20705 3565
rect 20725 3485 20735 3565
rect 20695 3475 20735 3485
<< mvpdiff >>
rect 9175 4305 9215 4315
rect 9175 4225 9185 4305
rect 9205 4225 9215 4305
rect 9175 4215 9215 4225
rect 9265 4305 9305 4315
rect 9265 4225 9275 4305
rect 9295 4225 9305 4305
rect 9265 4215 9305 4225
rect 9355 4305 9395 4315
rect 9355 4225 9365 4305
rect 9385 4225 9395 4305
rect 9355 4215 9395 4225
rect 9445 4305 9485 4315
rect 9445 4225 9455 4305
rect 9475 4225 9485 4305
rect 9445 4215 9485 4225
rect 9535 4305 9575 4315
rect 9535 4225 9545 4305
rect 9565 4225 9575 4305
rect 9535 4215 9575 4225
rect 9625 4305 9665 4315
rect 9625 4225 9635 4305
rect 9655 4225 9665 4305
rect 9625 4215 9665 4225
rect 9715 4305 9755 4315
rect 9715 4225 9725 4305
rect 9745 4225 9755 4305
rect 9715 4215 9755 4225
rect 9805 4305 9845 4315
rect 9805 4225 9815 4305
rect 9835 4225 9845 4305
rect 9805 4215 9845 4225
rect 9895 4305 9935 4315
rect 9895 4225 9905 4305
rect 9925 4225 9935 4305
rect 9895 4215 9935 4225
rect 9985 4305 10025 4315
rect 9985 4225 9995 4305
rect 10015 4225 10025 4305
rect 9985 4215 10025 4225
rect 10075 4305 10115 4315
rect 10075 4225 10085 4305
rect 10105 4225 10115 4305
rect 10075 4215 10115 4225
rect 10165 4305 10205 4315
rect 10165 4225 10175 4305
rect 10195 4225 10205 4305
rect 10165 4215 10205 4225
rect 10255 4305 10295 4315
rect 10255 4225 10265 4305
rect 10285 4225 10295 4305
rect 10255 4215 10295 4225
rect 10345 4305 10385 4315
rect 10345 4225 10355 4305
rect 10375 4225 10385 4305
rect 10345 4215 10385 4225
rect 10435 4305 10475 4315
rect 10435 4225 10445 4305
rect 10465 4225 10475 4305
rect 10435 4215 10475 4225
rect 10525 4305 10565 4315
rect 10525 4225 10535 4305
rect 10555 4225 10565 4305
rect 10525 4215 10565 4225
rect 10615 4305 10655 4315
rect 10615 4225 10625 4305
rect 10645 4225 10655 4305
rect 10615 4215 10655 4225
rect 10705 4305 10745 4315
rect 10705 4225 10715 4305
rect 10735 4225 10745 4305
rect 10705 4215 10745 4225
rect 10795 4305 10835 4315
rect 10795 4225 10805 4305
rect 10825 4225 10835 4305
rect 10795 4215 10835 4225
rect 10885 4305 10925 4315
rect 10885 4225 10895 4305
rect 10915 4225 10925 4305
rect 10885 4215 10925 4225
rect 10975 4305 11015 4315
rect 10975 4225 10985 4305
rect 11005 4225 11015 4305
rect 10975 4215 11015 4225
rect 11065 4305 11105 4315
rect 11065 4225 11075 4305
rect 11095 4225 11105 4305
rect 11065 4215 11105 4225
rect 11155 4305 11195 4315
rect 11155 4225 11165 4305
rect 11185 4225 11195 4305
rect 11155 4215 11195 4225
rect 11245 4305 11285 4315
rect 11245 4225 11255 4305
rect 11275 4225 11285 4305
rect 11245 4215 11285 4225
rect 11335 4305 11375 4315
rect 11335 4225 11345 4305
rect 11365 4225 11375 4305
rect 11335 4215 11375 4225
rect 11425 4305 11465 4315
rect 11425 4225 11435 4305
rect 11455 4225 11465 4305
rect 11425 4215 11465 4225
rect 11515 4305 11555 4315
rect 11515 4225 11525 4305
rect 11545 4225 11555 4305
rect 11515 4215 11555 4225
rect 11605 4305 11645 4315
rect 11605 4225 11615 4305
rect 11635 4225 11645 4305
rect 11605 4215 11645 4225
rect 11695 4305 11735 4315
rect 11695 4225 11705 4305
rect 11725 4225 11735 4305
rect 11695 4215 11735 4225
rect 11785 4305 11825 4315
rect 11785 4225 11795 4305
rect 11815 4225 11825 4305
rect 11785 4215 11825 4225
rect 11875 4305 11915 4315
rect 11875 4225 11885 4305
rect 11905 4225 11915 4305
rect 11875 4215 11915 4225
rect 11965 4305 12005 4315
rect 11965 4225 11975 4305
rect 11995 4225 12005 4305
rect 11965 4215 12005 4225
rect 12055 4305 12095 4315
rect 12055 4225 12065 4305
rect 12085 4225 12095 4305
rect 12055 4215 12095 4225
rect 12145 4305 12185 4315
rect 12145 4225 12155 4305
rect 12175 4225 12185 4305
rect 12145 4215 12185 4225
rect 12235 4305 12275 4315
rect 12235 4225 12245 4305
rect 12265 4225 12275 4305
rect 12235 4215 12275 4225
rect 12325 4305 12365 4315
rect 12325 4225 12335 4305
rect 12355 4225 12365 4305
rect 12325 4215 12365 4225
rect 12415 4305 12455 4315
rect 12415 4225 12425 4305
rect 12445 4225 12455 4305
rect 12415 4215 12455 4225
rect 12505 4305 12545 4315
rect 12505 4225 12515 4305
rect 12535 4225 12545 4305
rect 12505 4215 12545 4225
rect 12595 4305 12635 4315
rect 12595 4225 12605 4305
rect 12625 4225 12635 4305
rect 12595 4215 12635 4225
rect 12685 4305 12725 4315
rect 12685 4225 12695 4305
rect 12715 4225 12725 4305
rect 12685 4215 12725 4225
rect 12775 4305 12815 4315
rect 12775 4225 12785 4305
rect 12805 4225 12815 4305
rect 12775 4215 12815 4225
rect 12865 4305 12905 4315
rect 12865 4225 12875 4305
rect 12895 4225 12905 4305
rect 12865 4215 12905 4225
rect 12955 4305 12995 4315
rect 12955 4225 12965 4305
rect 12985 4225 12995 4305
rect 12955 4215 12995 4225
rect 13045 4305 13085 4315
rect 13045 4225 13055 4305
rect 13075 4225 13085 4305
rect 13045 4215 13085 4225
rect 13135 4305 13175 4315
rect 13135 4225 13145 4305
rect 13165 4225 13175 4305
rect 13135 4215 13175 4225
rect 13225 4305 13265 4315
rect 13225 4225 13235 4305
rect 13255 4225 13265 4305
rect 13225 4215 13265 4225
rect 13315 4305 13355 4315
rect 13315 4225 13325 4305
rect 13345 4225 13355 4305
rect 13315 4215 13355 4225
rect 13405 4305 13445 4315
rect 13405 4225 13415 4305
rect 13435 4225 13445 4305
rect 13405 4215 13445 4225
rect 13495 4305 13535 4315
rect 13495 4225 13505 4305
rect 13525 4225 13535 4305
rect 13495 4215 13535 4225
rect 13585 4305 13625 4315
rect 13585 4225 13595 4305
rect 13615 4225 13625 4305
rect 13585 4215 13625 4225
rect 13675 4305 13715 4315
rect 13675 4225 13685 4305
rect 13705 4225 13715 4305
rect 13675 4215 13715 4225
rect 13765 4305 13805 4315
rect 13765 4225 13775 4305
rect 13795 4225 13805 4305
rect 13765 4215 13805 4225
rect 13855 4305 13895 4315
rect 13855 4225 13865 4305
rect 13885 4225 13895 4305
rect 13855 4215 13895 4225
rect 13945 4305 13985 4315
rect 13945 4225 13955 4305
rect 13975 4225 13985 4305
rect 13945 4215 13985 4225
rect 14035 4305 14075 4315
rect 14035 4225 14045 4305
rect 14065 4225 14075 4305
rect 14035 4215 14075 4225
rect 14125 4305 14165 4315
rect 14125 4225 14135 4305
rect 14155 4225 14165 4305
rect 14125 4215 14165 4225
rect 14215 4305 14255 4315
rect 14215 4225 14225 4305
rect 14245 4225 14255 4305
rect 14215 4215 14255 4225
rect 14305 4305 14345 4315
rect 14305 4225 14315 4305
rect 14335 4225 14345 4305
rect 14305 4215 14345 4225
rect 14395 4305 14435 4315
rect 14395 4225 14405 4305
rect 14425 4225 14435 4305
rect 14395 4215 14435 4225
rect 14485 4305 14525 4315
rect 14485 4225 14495 4305
rect 14515 4225 14525 4305
rect 14485 4215 14525 4225
rect 14575 4305 14615 4315
rect 14575 4225 14585 4305
rect 14605 4225 14615 4305
rect 14575 4215 14615 4225
rect 14665 4305 14705 4315
rect 14665 4225 14675 4305
rect 14695 4225 14705 4305
rect 14665 4215 14705 4225
rect 14755 4305 14795 4315
rect 14755 4225 14765 4305
rect 14785 4225 14795 4305
rect 14755 4215 14795 4225
rect 14845 4305 14885 4315
rect 14845 4225 14855 4305
rect 14875 4225 14885 4305
rect 14845 4215 14885 4225
rect 14935 4305 14975 4315
rect 14935 4225 14945 4305
rect 14965 4225 14975 4305
rect 14935 4215 14975 4225
rect 15025 4305 15065 4315
rect 15025 4225 15035 4305
rect 15055 4225 15065 4305
rect 15025 4215 15065 4225
rect 15115 4305 15155 4315
rect 15115 4225 15125 4305
rect 15145 4225 15155 4305
rect 15115 4215 15155 4225
rect 15205 4305 15245 4315
rect 15205 4225 15215 4305
rect 15235 4225 15245 4305
rect 15205 4215 15245 4225
rect 15295 4305 15335 4315
rect 15295 4225 15305 4305
rect 15325 4225 15335 4305
rect 15295 4215 15335 4225
rect 15385 4305 15425 4315
rect 15385 4225 15395 4305
rect 15415 4225 15425 4305
rect 15385 4215 15425 4225
rect 15475 4305 15515 4315
rect 15475 4225 15485 4305
rect 15505 4225 15515 4305
rect 15475 4215 15515 4225
rect 15565 4305 15605 4315
rect 15565 4225 15575 4305
rect 15595 4225 15605 4305
rect 15565 4215 15605 4225
rect 15655 4305 15695 4315
rect 15655 4225 15665 4305
rect 15685 4225 15695 4305
rect 15655 4215 15695 4225
rect 15745 4305 15785 4315
rect 15745 4225 15755 4305
rect 15775 4225 15785 4305
rect 15745 4215 15785 4225
rect 15835 4305 15875 4315
rect 15835 4225 15845 4305
rect 15865 4225 15875 4305
rect 15835 4215 15875 4225
rect 15925 4305 15965 4315
rect 15925 4225 15935 4305
rect 15955 4225 15965 4305
rect 15925 4215 15965 4225
rect 16015 4305 16055 4315
rect 16015 4225 16025 4305
rect 16045 4225 16055 4305
rect 16015 4215 16055 4225
rect 16105 4305 16145 4315
rect 16105 4225 16115 4305
rect 16135 4225 16145 4305
rect 16105 4215 16145 4225
rect 16195 4305 16235 4315
rect 16195 4225 16205 4305
rect 16225 4225 16235 4305
rect 16195 4215 16235 4225
rect 16285 4305 16325 4315
rect 16285 4225 16295 4305
rect 16315 4225 16325 4305
rect 16285 4215 16325 4225
rect 16375 4305 16415 4315
rect 16375 4225 16385 4305
rect 16405 4225 16415 4305
rect 16375 4215 16415 4225
rect 16465 4305 16505 4315
rect 16465 4225 16475 4305
rect 16495 4225 16505 4305
rect 16465 4215 16505 4225
rect 16555 4305 16595 4315
rect 16555 4225 16565 4305
rect 16585 4225 16595 4305
rect 16555 4215 16595 4225
rect 16645 4305 16685 4315
rect 16645 4225 16655 4305
rect 16675 4225 16685 4305
rect 16645 4215 16685 4225
rect 16735 4305 16775 4315
rect 16735 4225 16745 4305
rect 16765 4225 16775 4305
rect 16735 4215 16775 4225
rect 16825 4305 16865 4315
rect 16825 4225 16835 4305
rect 16855 4225 16865 4305
rect 16825 4215 16865 4225
rect 16915 4305 16955 4315
rect 16915 4225 16925 4305
rect 16945 4225 16955 4305
rect 16915 4215 16955 4225
rect 17005 4305 17045 4315
rect 17005 4225 17015 4305
rect 17035 4225 17045 4305
rect 17005 4215 17045 4225
rect 17095 4305 17135 4315
rect 17095 4225 17105 4305
rect 17125 4225 17135 4305
rect 17095 4215 17135 4225
rect 17185 4305 17225 4315
rect 17185 4225 17195 4305
rect 17215 4225 17225 4305
rect 17185 4215 17225 4225
rect 17275 4305 17315 4315
rect 17275 4225 17285 4305
rect 17305 4225 17315 4305
rect 17275 4215 17315 4225
rect 17365 4305 17405 4315
rect 17365 4225 17375 4305
rect 17395 4225 17405 4305
rect 17365 4215 17405 4225
rect 17455 4305 17495 4315
rect 17455 4225 17465 4305
rect 17485 4225 17495 4305
rect 17455 4215 17495 4225
rect 17545 4305 17585 4315
rect 17545 4225 17555 4305
rect 17575 4225 17585 4305
rect 17545 4215 17585 4225
rect 17635 4305 17675 4315
rect 17635 4225 17645 4305
rect 17665 4225 17675 4305
rect 17635 4215 17675 4225
rect 17725 4305 17765 4315
rect 17725 4225 17735 4305
rect 17755 4225 17765 4305
rect 17725 4215 17765 4225
rect 17815 4305 17855 4315
rect 17815 4225 17825 4305
rect 17845 4225 17855 4305
rect 17815 4215 17855 4225
rect 17905 4305 17945 4315
rect 17905 4225 17915 4305
rect 17935 4225 17945 4305
rect 17905 4215 17945 4225
rect 17995 4305 18035 4315
rect 17995 4225 18005 4305
rect 18025 4225 18035 4305
rect 17995 4215 18035 4225
rect 18085 4305 18125 4315
rect 18085 4225 18095 4305
rect 18115 4225 18125 4305
rect 18085 4215 18125 4225
rect 18175 4305 18215 4315
rect 18175 4225 18185 4305
rect 18205 4225 18215 4305
rect 18175 4215 18215 4225
rect 18265 4305 18305 4315
rect 18265 4225 18275 4305
rect 18295 4225 18305 4305
rect 18265 4215 18305 4225
rect 18355 4305 18395 4315
rect 18355 4225 18365 4305
rect 18385 4225 18395 4305
rect 18355 4215 18395 4225
rect 18445 4305 18485 4315
rect 18445 4225 18455 4305
rect 18475 4225 18485 4305
rect 18445 4215 18485 4225
rect 18535 4305 18575 4315
rect 18535 4225 18545 4305
rect 18565 4225 18575 4305
rect 18535 4215 18575 4225
rect 18625 4305 18665 4315
rect 18625 4225 18635 4305
rect 18655 4225 18665 4305
rect 18625 4215 18665 4225
rect 18715 4305 18755 4315
rect 18715 4225 18725 4305
rect 18745 4225 18755 4305
rect 18715 4215 18755 4225
rect 18805 4305 18845 4315
rect 18805 4225 18815 4305
rect 18835 4225 18845 4305
rect 18805 4215 18845 4225
rect 18895 4305 18935 4315
rect 18895 4225 18905 4305
rect 18925 4225 18935 4305
rect 18895 4215 18935 4225
rect 18985 4305 19025 4315
rect 18985 4225 18995 4305
rect 19015 4225 19025 4305
rect 18985 4215 19025 4225
rect 19075 4305 19115 4315
rect 19075 4225 19085 4305
rect 19105 4225 19115 4305
rect 19075 4215 19115 4225
rect 19165 4305 19205 4315
rect 19165 4225 19175 4305
rect 19195 4225 19205 4305
rect 19165 4215 19205 4225
rect 19255 4305 19295 4315
rect 19255 4225 19265 4305
rect 19285 4225 19295 4305
rect 19255 4215 19295 4225
rect 19345 4305 19385 4315
rect 19345 4225 19355 4305
rect 19375 4225 19385 4305
rect 19345 4215 19385 4225
rect 19435 4305 19475 4315
rect 19435 4225 19445 4305
rect 19465 4225 19475 4305
rect 19435 4215 19475 4225
rect 19525 4305 19565 4315
rect 19525 4225 19535 4305
rect 19555 4225 19565 4305
rect 19525 4215 19565 4225
rect 19615 4305 19655 4315
rect 19615 4225 19625 4305
rect 19645 4225 19655 4305
rect 19615 4215 19655 4225
rect 19705 4305 19745 4315
rect 19705 4225 19715 4305
rect 19735 4225 19745 4305
rect 19705 4215 19745 4225
rect 19795 4305 19835 4315
rect 19795 4225 19805 4305
rect 19825 4225 19835 4305
rect 19795 4215 19835 4225
rect 19885 4305 19925 4315
rect 19885 4225 19895 4305
rect 19915 4225 19925 4305
rect 19885 4215 19925 4225
rect 19975 4305 20015 4315
rect 19975 4225 19985 4305
rect 20005 4225 20015 4305
rect 19975 4215 20015 4225
rect 20065 4305 20105 4315
rect 20065 4225 20075 4305
rect 20095 4225 20105 4305
rect 20065 4215 20105 4225
rect 20155 4305 20195 4315
rect 20155 4225 20165 4305
rect 20185 4225 20195 4305
rect 20155 4215 20195 4225
rect 20245 4305 20285 4315
rect 20245 4225 20255 4305
rect 20275 4225 20285 4305
rect 20245 4215 20285 4225
rect 20335 4305 20375 4315
rect 20335 4225 20345 4305
rect 20365 4225 20375 4305
rect 20335 4215 20375 4225
rect 20425 4305 20465 4315
rect 20425 4225 20435 4305
rect 20455 4225 20465 4305
rect 20425 4215 20465 4225
rect 20515 4305 20555 4315
rect 20515 4225 20525 4305
rect 20545 4225 20555 4305
rect 20515 4215 20555 4225
rect 20605 4305 20645 4315
rect 20605 4225 20615 4305
rect 20635 4225 20645 4305
rect 20605 4215 20645 4225
rect 20695 4305 20735 4315
rect 20695 4225 20705 4305
rect 20725 4225 20735 4305
rect 20695 4215 20735 4225
<< mvndiffc >>
rect 9185 3485 9205 3565
rect 9275 3485 9295 3565
rect 9365 3485 9385 3565
rect 9455 3485 9475 3565
rect 9545 3485 9565 3565
rect 9635 3485 9655 3565
rect 9725 3485 9745 3565
rect 9815 3485 9835 3565
rect 9905 3485 9925 3565
rect 9995 3485 10015 3565
rect 10085 3485 10105 3565
rect 10175 3485 10195 3565
rect 10265 3485 10285 3565
rect 10355 3485 10375 3565
rect 10445 3485 10465 3565
rect 10535 3485 10555 3565
rect 10625 3485 10645 3565
rect 10715 3485 10735 3565
rect 10805 3485 10825 3565
rect 10895 3485 10915 3565
rect 10985 3485 11005 3565
rect 11075 3485 11095 3565
rect 11165 3485 11185 3565
rect 11255 3485 11275 3565
rect 11345 3485 11365 3565
rect 11435 3485 11455 3565
rect 11525 3485 11545 3565
rect 11615 3485 11635 3565
rect 11705 3485 11725 3565
rect 11795 3485 11815 3565
rect 11885 3485 11905 3565
rect 11975 3485 11995 3565
rect 12065 3485 12085 3565
rect 12155 3485 12175 3565
rect 12245 3485 12265 3565
rect 12335 3485 12355 3565
rect 12425 3485 12445 3565
rect 12515 3485 12535 3565
rect 12605 3485 12625 3565
rect 12695 3485 12715 3565
rect 12785 3485 12805 3565
rect 12875 3485 12895 3565
rect 12965 3485 12985 3565
rect 13055 3485 13075 3565
rect 13145 3485 13165 3565
rect 13235 3485 13255 3565
rect 13325 3485 13345 3565
rect 13415 3485 13435 3565
rect 13505 3485 13525 3565
rect 13595 3485 13615 3565
rect 13685 3485 13705 3565
rect 13775 3485 13795 3565
rect 13865 3485 13885 3565
rect 13955 3485 13975 3565
rect 14045 3485 14065 3565
rect 14135 3485 14155 3565
rect 14225 3485 14245 3565
rect 14315 3485 14335 3565
rect 14405 3485 14425 3565
rect 14495 3485 14515 3565
rect 14585 3485 14605 3565
rect 14675 3485 14695 3565
rect 14765 3485 14785 3565
rect 14855 3485 14875 3565
rect 14945 3485 14965 3565
rect 15035 3485 15055 3565
rect 15125 3485 15145 3565
rect 15215 3485 15235 3565
rect 15305 3485 15325 3565
rect 15395 3485 15415 3565
rect 15485 3485 15505 3565
rect 15575 3485 15595 3565
rect 15665 3485 15685 3565
rect 15755 3485 15775 3565
rect 15845 3485 15865 3565
rect 15935 3485 15955 3565
rect 16025 3485 16045 3565
rect 16115 3485 16135 3565
rect 16205 3485 16225 3565
rect 16295 3485 16315 3565
rect 16385 3485 16405 3565
rect 16475 3485 16495 3565
rect 16565 3485 16585 3565
rect 16655 3485 16675 3565
rect 16745 3485 16765 3565
rect 16835 3485 16855 3565
rect 16925 3485 16945 3565
rect 17015 3485 17035 3565
rect 17105 3485 17125 3565
rect 17195 3485 17215 3565
rect 17285 3485 17305 3565
rect 17375 3485 17395 3565
rect 17465 3485 17485 3565
rect 17555 3485 17575 3565
rect 17645 3485 17665 3565
rect 17735 3485 17755 3565
rect 17825 3485 17845 3565
rect 17915 3485 17935 3565
rect 18005 3485 18025 3565
rect 18095 3485 18115 3565
rect 18185 3485 18205 3565
rect 18275 3485 18295 3565
rect 18365 3485 18385 3565
rect 18455 3485 18475 3565
rect 18545 3485 18565 3565
rect 18635 3485 18655 3565
rect 18725 3485 18745 3565
rect 18815 3485 18835 3565
rect 18905 3485 18925 3565
rect 18995 3485 19015 3565
rect 19085 3485 19105 3565
rect 19175 3485 19195 3565
rect 19265 3485 19285 3565
rect 19355 3485 19375 3565
rect 19445 3485 19465 3565
rect 19535 3485 19555 3565
rect 19625 3485 19645 3565
rect 19715 3485 19735 3565
rect 19805 3485 19825 3565
rect 19895 3485 19915 3565
rect 19985 3485 20005 3565
rect 20075 3485 20095 3565
rect 20165 3485 20185 3565
rect 20255 3485 20275 3565
rect 20345 3485 20365 3565
rect 20435 3485 20455 3565
rect 20525 3485 20545 3565
rect 20615 3485 20635 3565
rect 20705 3485 20725 3565
<< mvpdiffc >>
rect 9185 4225 9205 4305
rect 9275 4225 9295 4305
rect 9365 4225 9385 4305
rect 9455 4225 9475 4305
rect 9545 4225 9565 4305
rect 9635 4225 9655 4305
rect 9725 4225 9745 4305
rect 9815 4225 9835 4305
rect 9905 4225 9925 4305
rect 9995 4225 10015 4305
rect 10085 4225 10105 4305
rect 10175 4225 10195 4305
rect 10265 4225 10285 4305
rect 10355 4225 10375 4305
rect 10445 4225 10465 4305
rect 10535 4225 10555 4305
rect 10625 4225 10645 4305
rect 10715 4225 10735 4305
rect 10805 4225 10825 4305
rect 10895 4225 10915 4305
rect 10985 4225 11005 4305
rect 11075 4225 11095 4305
rect 11165 4225 11185 4305
rect 11255 4225 11275 4305
rect 11345 4225 11365 4305
rect 11435 4225 11455 4305
rect 11525 4225 11545 4305
rect 11615 4225 11635 4305
rect 11705 4225 11725 4305
rect 11795 4225 11815 4305
rect 11885 4225 11905 4305
rect 11975 4225 11995 4305
rect 12065 4225 12085 4305
rect 12155 4225 12175 4305
rect 12245 4225 12265 4305
rect 12335 4225 12355 4305
rect 12425 4225 12445 4305
rect 12515 4225 12535 4305
rect 12605 4225 12625 4305
rect 12695 4225 12715 4305
rect 12785 4225 12805 4305
rect 12875 4225 12895 4305
rect 12965 4225 12985 4305
rect 13055 4225 13075 4305
rect 13145 4225 13165 4305
rect 13235 4225 13255 4305
rect 13325 4225 13345 4305
rect 13415 4225 13435 4305
rect 13505 4225 13525 4305
rect 13595 4225 13615 4305
rect 13685 4225 13705 4305
rect 13775 4225 13795 4305
rect 13865 4225 13885 4305
rect 13955 4225 13975 4305
rect 14045 4225 14065 4305
rect 14135 4225 14155 4305
rect 14225 4225 14245 4305
rect 14315 4225 14335 4305
rect 14405 4225 14425 4305
rect 14495 4225 14515 4305
rect 14585 4225 14605 4305
rect 14675 4225 14695 4305
rect 14765 4225 14785 4305
rect 14855 4225 14875 4305
rect 14945 4225 14965 4305
rect 15035 4225 15055 4305
rect 15125 4225 15145 4305
rect 15215 4225 15235 4305
rect 15305 4225 15325 4305
rect 15395 4225 15415 4305
rect 15485 4225 15505 4305
rect 15575 4225 15595 4305
rect 15665 4225 15685 4305
rect 15755 4225 15775 4305
rect 15845 4225 15865 4305
rect 15935 4225 15955 4305
rect 16025 4225 16045 4305
rect 16115 4225 16135 4305
rect 16205 4225 16225 4305
rect 16295 4225 16315 4305
rect 16385 4225 16405 4305
rect 16475 4225 16495 4305
rect 16565 4225 16585 4305
rect 16655 4225 16675 4305
rect 16745 4225 16765 4305
rect 16835 4225 16855 4305
rect 16925 4225 16945 4305
rect 17015 4225 17035 4305
rect 17105 4225 17125 4305
rect 17195 4225 17215 4305
rect 17285 4225 17305 4305
rect 17375 4225 17395 4305
rect 17465 4225 17485 4305
rect 17555 4225 17575 4305
rect 17645 4225 17665 4305
rect 17735 4225 17755 4305
rect 17825 4225 17845 4305
rect 17915 4225 17935 4305
rect 18005 4225 18025 4305
rect 18095 4225 18115 4305
rect 18185 4225 18205 4305
rect 18275 4225 18295 4305
rect 18365 4225 18385 4305
rect 18455 4225 18475 4305
rect 18545 4225 18565 4305
rect 18635 4225 18655 4305
rect 18725 4225 18745 4305
rect 18815 4225 18835 4305
rect 18905 4225 18925 4305
rect 18995 4225 19015 4305
rect 19085 4225 19105 4305
rect 19175 4225 19195 4305
rect 19265 4225 19285 4305
rect 19355 4225 19375 4305
rect 19445 4225 19465 4305
rect 19535 4225 19555 4305
rect 19625 4225 19645 4305
rect 19715 4225 19735 4305
rect 19805 4225 19825 4305
rect 19895 4225 19915 4305
rect 19985 4225 20005 4305
rect 20075 4225 20095 4305
rect 20165 4225 20185 4305
rect 20255 4225 20275 4305
rect 20345 4225 20365 4305
rect 20435 4225 20455 4305
rect 20525 4225 20545 4305
rect 20615 4225 20635 4305
rect 20705 4225 20725 4305
<< psubdiff >>
rect 9050 4065 9070 4375
rect 20840 4065 20860 4375
rect 9050 4045 9230 4065
rect 9250 4045 9320 4065
rect 9340 4045 9410 4065
rect 9430 4045 9500 4065
rect 9520 4045 9590 4065
rect 9610 4045 9680 4065
rect 9700 4045 9770 4065
rect 9790 4045 9860 4065
rect 9880 4045 9950 4065
rect 9970 4045 10040 4065
rect 10060 4045 10130 4065
rect 10150 4045 10220 4065
rect 10240 4045 10310 4065
rect 10330 4045 10400 4065
rect 10420 4045 10490 4065
rect 10510 4045 10580 4065
rect 10600 4045 10670 4065
rect 10690 4045 10760 4065
rect 10780 4045 10850 4065
rect 10870 4045 10940 4065
rect 10960 4045 11030 4065
rect 11050 4045 11120 4065
rect 11140 4045 11210 4065
rect 11230 4045 11300 4065
rect 11320 4045 11390 4065
rect 11410 4045 11480 4065
rect 11500 4045 11570 4065
rect 11590 4045 11660 4065
rect 11680 4045 11750 4065
rect 11770 4045 11840 4065
rect 11860 4045 11930 4065
rect 11950 4045 12020 4065
rect 12040 4045 12110 4065
rect 12130 4045 12200 4065
rect 12220 4045 12290 4065
rect 12310 4045 12380 4065
rect 12400 4045 12470 4065
rect 12490 4045 12560 4065
rect 12580 4045 12650 4065
rect 12670 4045 12740 4065
rect 12760 4045 12830 4065
rect 12850 4045 12920 4065
rect 12940 4045 13010 4065
rect 13030 4045 13100 4065
rect 13120 4045 13190 4065
rect 13210 4045 13280 4065
rect 13300 4045 13370 4065
rect 13390 4045 13460 4065
rect 13480 4045 13550 4065
rect 13570 4045 13640 4065
rect 13660 4045 13730 4065
rect 13750 4045 13820 4065
rect 13840 4045 13910 4065
rect 13930 4045 14000 4065
rect 14020 4045 14090 4065
rect 14110 4045 14180 4065
rect 14200 4045 14270 4065
rect 14290 4045 14360 4065
rect 14380 4045 14450 4065
rect 14470 4045 14540 4065
rect 14560 4045 14630 4065
rect 14650 4045 14720 4065
rect 14740 4045 14810 4065
rect 14830 4045 14900 4065
rect 14920 4045 14990 4065
rect 15010 4045 15080 4065
rect 15100 4045 15170 4065
rect 15190 4045 15260 4065
rect 15280 4045 15350 4065
rect 15370 4045 15440 4065
rect 15460 4045 15530 4065
rect 15550 4045 15620 4065
rect 15640 4045 15710 4065
rect 15730 4045 15800 4065
rect 15820 4045 15890 4065
rect 15910 4045 15980 4065
rect 16000 4045 16070 4065
rect 16090 4045 16160 4065
rect 16180 4045 16250 4065
rect 16270 4045 16340 4065
rect 16360 4045 16430 4065
rect 16450 4045 16520 4065
rect 16540 4045 16610 4065
rect 16630 4045 16700 4065
rect 16720 4045 16790 4065
rect 16810 4045 16880 4065
rect 16900 4045 16970 4065
rect 16990 4045 17060 4065
rect 17080 4045 17150 4065
rect 17170 4045 17240 4065
rect 17260 4045 17330 4065
rect 17350 4045 17420 4065
rect 17440 4045 17510 4065
rect 17530 4045 17600 4065
rect 17620 4045 17690 4065
rect 17710 4045 17780 4065
rect 17800 4045 17870 4065
rect 17890 4045 17960 4065
rect 17980 4045 18050 4065
rect 18070 4045 18140 4065
rect 18160 4045 18230 4065
rect 18250 4045 18320 4065
rect 18340 4045 18410 4065
rect 18430 4045 18500 4065
rect 18520 4045 18590 4065
rect 18610 4045 18680 4065
rect 18700 4045 18770 4065
rect 18790 4045 18860 4065
rect 18880 4045 18950 4065
rect 18970 4045 19040 4065
rect 19060 4045 19130 4065
rect 19150 4045 19220 4065
rect 19240 4045 19310 4065
rect 19330 4045 19400 4065
rect 19420 4045 19490 4065
rect 19510 4045 19580 4065
rect 19600 4045 19670 4065
rect 19690 4045 19760 4065
rect 19780 4045 19850 4065
rect 19870 4045 19940 4065
rect 19960 4045 20030 4065
rect 20050 4045 20120 4065
rect 20140 4045 20210 4065
rect 20230 4045 20300 4065
rect 20320 4045 20390 4065
rect 20410 4045 20480 4065
rect 20500 4045 20570 4065
rect 20590 4045 20660 4065
rect 20680 4045 20860 4065
rect 9050 3645 9230 3665
rect 9250 3645 9320 3665
rect 9340 3645 9410 3665
rect 9430 3645 9500 3665
rect 9520 3645 9590 3665
rect 9610 3645 9680 3665
rect 9700 3645 9770 3665
rect 9790 3645 9860 3665
rect 9880 3645 9950 3665
rect 9970 3645 10040 3665
rect 10060 3645 10130 3665
rect 10150 3645 10220 3665
rect 10240 3645 10310 3665
rect 10330 3645 10400 3665
rect 10420 3645 10490 3665
rect 10510 3645 10580 3665
rect 10600 3645 10670 3665
rect 10690 3645 10760 3665
rect 10780 3645 10850 3665
rect 10870 3645 10940 3665
rect 10960 3645 11030 3665
rect 11050 3645 11120 3665
rect 11140 3645 11210 3665
rect 11230 3645 11300 3665
rect 11320 3645 11390 3665
rect 11410 3645 11480 3665
rect 11500 3645 11570 3665
rect 11590 3645 11660 3665
rect 11680 3645 11750 3665
rect 11770 3645 11840 3665
rect 11860 3645 11930 3665
rect 11950 3645 12020 3665
rect 12040 3645 12110 3665
rect 12130 3645 12200 3665
rect 12220 3645 12290 3665
rect 12310 3645 12380 3665
rect 12400 3645 12470 3665
rect 12490 3645 12560 3665
rect 12580 3645 12650 3665
rect 12670 3645 12740 3665
rect 12760 3645 12830 3665
rect 12850 3645 12920 3665
rect 12940 3645 13010 3665
rect 13030 3645 13100 3665
rect 13120 3645 13190 3665
rect 13210 3645 13280 3665
rect 13300 3645 13370 3665
rect 13390 3645 13460 3665
rect 13480 3645 13550 3665
rect 13570 3645 13640 3665
rect 13660 3645 13730 3665
rect 13750 3645 13820 3665
rect 13840 3645 13910 3665
rect 13930 3645 14000 3665
rect 14020 3645 14090 3665
rect 14110 3645 14180 3665
rect 14200 3645 14270 3665
rect 14290 3645 14360 3665
rect 14380 3645 14450 3665
rect 14470 3645 14540 3665
rect 14560 3645 14630 3665
rect 14650 3645 14720 3665
rect 14740 3645 14810 3665
rect 14830 3645 14900 3665
rect 14920 3645 14990 3665
rect 15010 3645 15080 3665
rect 15100 3645 15170 3665
rect 15190 3645 15260 3665
rect 15280 3645 15350 3665
rect 15370 3645 15440 3665
rect 15460 3645 15530 3665
rect 15550 3645 15620 3665
rect 15640 3645 15710 3665
rect 15730 3645 15800 3665
rect 15820 3645 15890 3665
rect 15910 3645 15980 3665
rect 16000 3645 16070 3665
rect 16090 3645 16160 3665
rect 16180 3645 16250 3665
rect 16270 3645 16340 3665
rect 16360 3645 16430 3665
rect 16450 3645 16520 3665
rect 16540 3645 16610 3665
rect 16630 3645 16700 3665
rect 16720 3645 16790 3665
rect 16810 3645 16880 3665
rect 16900 3645 16970 3665
rect 16990 3645 17060 3665
rect 17080 3645 17150 3665
rect 17170 3645 17240 3665
rect 17260 3645 17330 3665
rect 17350 3645 17420 3665
rect 17440 3645 17510 3665
rect 17530 3645 17600 3665
rect 17620 3645 17690 3665
rect 17710 3645 17780 3665
rect 17800 3645 17870 3665
rect 17890 3645 17960 3665
rect 17980 3645 18050 3665
rect 18070 3645 18140 3665
rect 18160 3645 18230 3665
rect 18250 3645 18320 3665
rect 18340 3645 18410 3665
rect 18430 3645 18500 3665
rect 18520 3645 18590 3665
rect 18610 3645 18680 3665
rect 18700 3645 18770 3665
rect 18790 3645 18860 3665
rect 18880 3645 18950 3665
rect 18970 3645 19040 3665
rect 19060 3645 19130 3665
rect 19150 3645 19220 3665
rect 19240 3645 19310 3665
rect 19330 3645 19400 3665
rect 19420 3645 19490 3665
rect 19510 3645 19580 3665
rect 19600 3645 19670 3665
rect 19690 3645 19760 3665
rect 19780 3645 19850 3665
rect 19870 3645 19940 3665
rect 19960 3645 20030 3665
rect 20050 3645 20120 3665
rect 20140 3645 20210 3665
rect 20230 3645 20300 3665
rect 20320 3645 20390 3665
rect 20410 3645 20480 3665
rect 20500 3645 20570 3665
rect 20590 3645 20660 3665
rect 20680 3645 20860 3665
rect 9050 3445 9070 3645
rect 20840 3445 20860 3645
rect 9040 3425 9230 3445
rect 9250 3425 9320 3445
rect 9340 3425 9410 3445
rect 9430 3425 9500 3445
rect 9520 3425 9590 3445
rect 9610 3425 9680 3445
rect 9700 3425 9770 3445
rect 9790 3425 9860 3445
rect 9880 3425 9950 3445
rect 9970 3425 10040 3445
rect 10060 3425 10130 3445
rect 10150 3425 10220 3445
rect 10240 3425 10310 3445
rect 10330 3425 10400 3445
rect 10420 3425 10490 3445
rect 10510 3425 10580 3445
rect 10600 3425 10670 3445
rect 10690 3425 10760 3445
rect 10780 3425 10850 3445
rect 10870 3425 10940 3445
rect 10960 3425 11030 3445
rect 11050 3425 11120 3445
rect 11140 3425 11210 3445
rect 11230 3425 11300 3445
rect 11320 3425 11390 3445
rect 11410 3425 11480 3445
rect 11500 3425 11570 3445
rect 11590 3425 11660 3445
rect 11680 3425 11750 3445
rect 11770 3425 11840 3445
rect 11860 3425 11930 3445
rect 11950 3425 12020 3445
rect 12040 3425 12110 3445
rect 12130 3425 12200 3445
rect 12220 3425 12290 3445
rect 12310 3425 12380 3445
rect 12400 3425 12470 3445
rect 12490 3425 12560 3445
rect 12580 3425 12650 3445
rect 12670 3425 12740 3445
rect 12760 3425 12830 3445
rect 12850 3425 12920 3445
rect 12940 3425 13010 3445
rect 13030 3425 13100 3445
rect 13120 3425 13190 3445
rect 13210 3425 13280 3445
rect 13300 3425 13370 3445
rect 13390 3425 13460 3445
rect 13480 3425 13550 3445
rect 13570 3425 13640 3445
rect 13660 3425 13730 3445
rect 13750 3425 13820 3445
rect 13840 3425 13910 3445
rect 13930 3425 14000 3445
rect 14020 3425 14090 3445
rect 14110 3425 14180 3445
rect 14200 3425 14270 3445
rect 14290 3425 14360 3445
rect 14380 3425 14450 3445
rect 14470 3425 14540 3445
rect 14560 3425 14630 3445
rect 14650 3425 14720 3445
rect 14740 3425 14810 3445
rect 14830 3425 14900 3445
rect 14920 3425 14990 3445
rect 15010 3425 15080 3445
rect 15100 3425 15170 3445
rect 15190 3425 15260 3445
rect 15280 3425 15350 3445
rect 15370 3425 15440 3445
rect 15460 3425 15530 3445
rect 15550 3425 15620 3445
rect 15640 3425 15710 3445
rect 15730 3425 15800 3445
rect 15820 3425 15890 3445
rect 15910 3425 15980 3445
rect 16000 3425 16070 3445
rect 16090 3425 16160 3445
rect 16180 3425 16250 3445
rect 16270 3425 16340 3445
rect 16360 3425 16430 3445
rect 16450 3425 16520 3445
rect 16540 3425 16610 3445
rect 16630 3425 16700 3445
rect 16720 3425 16790 3445
rect 16810 3425 16880 3445
rect 16900 3425 16970 3445
rect 16990 3425 17060 3445
rect 17080 3425 17150 3445
rect 17170 3425 17240 3445
rect 17260 3425 17330 3445
rect 17350 3425 17420 3445
rect 17440 3425 17510 3445
rect 17530 3425 17600 3445
rect 17620 3425 17690 3445
rect 17710 3425 17780 3445
rect 17800 3425 17870 3445
rect 17890 3425 17960 3445
rect 17980 3425 18050 3445
rect 18070 3425 18140 3445
rect 18160 3425 18230 3445
rect 18250 3425 18320 3445
rect 18340 3425 18410 3445
rect 18430 3425 18500 3445
rect 18520 3425 18590 3445
rect 18610 3425 18680 3445
rect 18700 3425 18770 3445
rect 18790 3425 18860 3445
rect 18880 3425 18950 3445
rect 18970 3425 19040 3445
rect 19060 3425 19130 3445
rect 19150 3425 19220 3445
rect 19240 3425 19310 3445
rect 19330 3425 19400 3445
rect 19420 3425 19490 3445
rect 19510 3425 19580 3445
rect 19600 3425 19670 3445
rect 19690 3425 19760 3445
rect 19780 3425 19850 3445
rect 19870 3425 19940 3445
rect 19960 3425 20030 3445
rect 20050 3425 20120 3445
rect 20140 3425 20210 3445
rect 20230 3425 20300 3445
rect 20320 3425 20390 3445
rect 20410 3425 20480 3445
rect 20500 3425 20570 3445
rect 20590 3425 20660 3445
rect 20680 3425 20870 3445
<< nsubdiff >>
rect 9125 4345 9230 4365
rect 9250 4345 9320 4365
rect 9340 4345 9410 4365
rect 9430 4345 9500 4365
rect 9520 4345 9590 4365
rect 9610 4345 9680 4365
rect 9700 4345 9770 4365
rect 9790 4345 9860 4365
rect 9880 4345 9950 4365
rect 9970 4345 10040 4365
rect 10060 4345 10130 4365
rect 10150 4345 10220 4365
rect 10240 4345 10310 4365
rect 10330 4345 10400 4365
rect 10420 4345 10490 4365
rect 10510 4345 10580 4365
rect 10600 4345 10670 4365
rect 10690 4345 10760 4365
rect 10780 4345 10850 4365
rect 10870 4345 10940 4365
rect 10960 4345 11030 4365
rect 11050 4345 11120 4365
rect 11140 4345 11210 4365
rect 11230 4345 11300 4365
rect 11320 4345 11390 4365
rect 11410 4345 11480 4365
rect 11500 4345 11570 4365
rect 11590 4345 11660 4365
rect 11680 4345 11750 4365
rect 11770 4345 11840 4365
rect 11860 4345 11930 4365
rect 11950 4345 12020 4365
rect 12040 4345 12110 4365
rect 12130 4345 12200 4365
rect 12220 4345 12290 4365
rect 12310 4345 12380 4365
rect 12400 4345 12470 4365
rect 12490 4345 12560 4365
rect 12580 4345 12650 4365
rect 12670 4345 12740 4365
rect 12760 4345 12830 4365
rect 12850 4345 12920 4365
rect 12940 4345 13010 4365
rect 13030 4345 13100 4365
rect 13120 4345 13190 4365
rect 13210 4345 13280 4365
rect 13300 4345 13370 4365
rect 13390 4345 13460 4365
rect 13480 4345 13550 4365
rect 13570 4345 13640 4365
rect 13660 4345 13730 4365
rect 13750 4345 13820 4365
rect 13840 4345 13910 4365
rect 13930 4345 14000 4365
rect 14020 4345 14090 4365
rect 14110 4345 14180 4365
rect 14200 4345 14270 4365
rect 14290 4345 14360 4365
rect 14380 4345 14450 4365
rect 14470 4345 14540 4365
rect 14560 4345 14630 4365
rect 14650 4345 14720 4365
rect 14740 4345 14810 4365
rect 14830 4345 14900 4365
rect 14920 4345 14990 4365
rect 15010 4345 15080 4365
rect 15100 4345 15170 4365
rect 15190 4345 15260 4365
rect 15280 4345 15350 4365
rect 15370 4345 15440 4365
rect 15460 4345 15530 4365
rect 15550 4345 15620 4365
rect 15640 4345 15710 4365
rect 15730 4345 15800 4365
rect 15820 4345 15890 4365
rect 15910 4345 15980 4365
rect 16000 4345 16070 4365
rect 16090 4345 16160 4365
rect 16180 4345 16250 4365
rect 16270 4345 16340 4365
rect 16360 4345 16430 4365
rect 16450 4345 16520 4365
rect 16540 4345 16610 4365
rect 16630 4345 16700 4365
rect 16720 4345 16790 4365
rect 16810 4345 16880 4365
rect 16900 4345 16970 4365
rect 16990 4345 17060 4365
rect 17080 4345 17150 4365
rect 17170 4345 17240 4365
rect 17260 4345 17330 4365
rect 17350 4345 17420 4365
rect 17440 4345 17510 4365
rect 17530 4345 17600 4365
rect 17620 4345 17690 4365
rect 17710 4345 17780 4365
rect 17800 4345 17870 4365
rect 17890 4345 17960 4365
rect 17980 4345 18050 4365
rect 18070 4345 18140 4365
rect 18160 4345 18230 4365
rect 18250 4345 18320 4365
rect 18340 4345 18410 4365
rect 18430 4345 18500 4365
rect 18520 4345 18590 4365
rect 18610 4345 18680 4365
rect 18700 4345 18770 4365
rect 18790 4345 18860 4365
rect 18880 4345 18950 4365
rect 18970 4345 19040 4365
rect 19060 4345 19130 4365
rect 19150 4345 19220 4365
rect 19240 4345 19310 4365
rect 19330 4345 19400 4365
rect 19420 4345 19490 4365
rect 19510 4345 19580 4365
rect 19600 4345 19670 4365
rect 19690 4345 19760 4365
rect 19780 4345 19850 4365
rect 19870 4345 19940 4365
rect 19960 4345 20030 4365
rect 20050 4345 20120 4365
rect 20140 4345 20210 4365
rect 20230 4345 20300 4365
rect 20320 4345 20390 4365
rect 20410 4345 20480 4365
rect 20500 4345 20570 4365
rect 20590 4345 20660 4365
rect 20680 4345 20785 4365
rect 9125 4145 9145 4345
rect 20765 4145 20785 4345
rect 9125 4125 9230 4145
rect 9250 4125 9320 4145
rect 9340 4125 9410 4145
rect 9430 4125 9500 4145
rect 9520 4125 9590 4145
rect 9610 4125 9680 4145
rect 9700 4125 9770 4145
rect 9790 4125 9860 4145
rect 9880 4125 9950 4145
rect 9970 4125 10040 4145
rect 10060 4125 10130 4145
rect 10150 4125 10220 4145
rect 10240 4125 10310 4145
rect 10330 4125 10400 4145
rect 10420 4125 10490 4145
rect 10510 4125 10580 4145
rect 10600 4125 10670 4145
rect 10690 4125 10760 4145
rect 10780 4125 10850 4145
rect 10870 4125 10940 4145
rect 10960 4125 11030 4145
rect 11050 4125 11120 4145
rect 11140 4125 11210 4145
rect 11230 4125 11300 4145
rect 11320 4125 11390 4145
rect 11410 4125 11480 4145
rect 11500 4125 11570 4145
rect 11590 4125 11660 4145
rect 11680 4125 11750 4145
rect 11770 4125 11840 4145
rect 11860 4125 11930 4145
rect 11950 4125 12020 4145
rect 12040 4125 12110 4145
rect 12130 4125 12200 4145
rect 12220 4125 12290 4145
rect 12310 4125 12380 4145
rect 12400 4125 12470 4145
rect 12490 4125 12560 4145
rect 12580 4125 12650 4145
rect 12670 4125 12740 4145
rect 12760 4125 12830 4145
rect 12850 4125 12920 4145
rect 12940 4125 13010 4145
rect 13030 4125 13100 4145
rect 13120 4125 13190 4145
rect 13210 4125 13280 4145
rect 13300 4125 13370 4145
rect 13390 4125 13460 4145
rect 13480 4125 13550 4145
rect 13570 4125 13640 4145
rect 13660 4125 13730 4145
rect 13750 4125 13820 4145
rect 13840 4125 13910 4145
rect 13930 4125 14000 4145
rect 14020 4125 14090 4145
rect 14110 4125 14180 4145
rect 14200 4125 14270 4145
rect 14290 4125 14360 4145
rect 14380 4125 14450 4145
rect 14470 4125 14540 4145
rect 14560 4125 14630 4145
rect 14650 4125 14720 4145
rect 14740 4125 14810 4145
rect 14830 4125 14900 4145
rect 14920 4125 14990 4145
rect 15010 4125 15080 4145
rect 15100 4125 15170 4145
rect 15190 4125 15260 4145
rect 15280 4125 15350 4145
rect 15370 4125 15440 4145
rect 15460 4125 15530 4145
rect 15550 4125 15620 4145
rect 15640 4125 15710 4145
rect 15730 4125 15800 4145
rect 15820 4125 15890 4145
rect 15910 4125 15980 4145
rect 16000 4125 16070 4145
rect 16090 4125 16160 4145
rect 16180 4125 16250 4145
rect 16270 4125 16340 4145
rect 16360 4125 16430 4145
rect 16450 4125 16520 4145
rect 16540 4125 16610 4145
rect 16630 4125 16700 4145
rect 16720 4125 16790 4145
rect 16810 4125 16880 4145
rect 16900 4125 16970 4145
rect 16990 4125 17060 4145
rect 17080 4125 17150 4145
rect 17170 4125 17240 4145
rect 17260 4125 17330 4145
rect 17350 4125 17420 4145
rect 17440 4125 17510 4145
rect 17530 4125 17600 4145
rect 17620 4125 17690 4145
rect 17710 4125 17780 4145
rect 17800 4125 17870 4145
rect 17890 4125 17960 4145
rect 17980 4125 18050 4145
rect 18070 4125 18140 4145
rect 18160 4125 18230 4145
rect 18250 4125 18320 4145
rect 18340 4125 18410 4145
rect 18430 4125 18500 4145
rect 18520 4125 18590 4145
rect 18610 4125 18680 4145
rect 18700 4125 18770 4145
rect 18790 4125 18860 4145
rect 18880 4125 18950 4145
rect 18970 4125 19040 4145
rect 19060 4125 19130 4145
rect 19150 4125 19220 4145
rect 19240 4125 19310 4145
rect 19330 4125 19400 4145
rect 19420 4125 19490 4145
rect 19510 4125 19580 4145
rect 19600 4125 19670 4145
rect 19690 4125 19760 4145
rect 19780 4125 19850 4145
rect 19870 4125 19940 4145
rect 19960 4125 20030 4145
rect 20050 4125 20120 4145
rect 20140 4125 20210 4145
rect 20230 4125 20300 4145
rect 20320 4125 20390 4145
rect 20410 4125 20480 4145
rect 20500 4125 20570 4145
rect 20590 4125 20660 4145
rect 20680 4125 20785 4145
<< psubdiffcont >>
rect 9230 4045 9250 4065
rect 9320 4045 9340 4065
rect 9410 4045 9430 4065
rect 9500 4045 9520 4065
rect 9590 4045 9610 4065
rect 9680 4045 9700 4065
rect 9770 4045 9790 4065
rect 9860 4045 9880 4065
rect 9950 4045 9970 4065
rect 10040 4045 10060 4065
rect 10130 4045 10150 4065
rect 10220 4045 10240 4065
rect 10310 4045 10330 4065
rect 10400 4045 10420 4065
rect 10490 4045 10510 4065
rect 10580 4045 10600 4065
rect 10670 4045 10690 4065
rect 10760 4045 10780 4065
rect 10850 4045 10870 4065
rect 10940 4045 10960 4065
rect 11030 4045 11050 4065
rect 11120 4045 11140 4065
rect 11210 4045 11230 4065
rect 11300 4045 11320 4065
rect 11390 4045 11410 4065
rect 11480 4045 11500 4065
rect 11570 4045 11590 4065
rect 11660 4045 11680 4065
rect 11750 4045 11770 4065
rect 11840 4045 11860 4065
rect 11930 4045 11950 4065
rect 12020 4045 12040 4065
rect 12110 4045 12130 4065
rect 12200 4045 12220 4065
rect 12290 4045 12310 4065
rect 12380 4045 12400 4065
rect 12470 4045 12490 4065
rect 12560 4045 12580 4065
rect 12650 4045 12670 4065
rect 12740 4045 12760 4065
rect 12830 4045 12850 4065
rect 12920 4045 12940 4065
rect 13010 4045 13030 4065
rect 13100 4045 13120 4065
rect 13190 4045 13210 4065
rect 13280 4045 13300 4065
rect 13370 4045 13390 4065
rect 13460 4045 13480 4065
rect 13550 4045 13570 4065
rect 13640 4045 13660 4065
rect 13730 4045 13750 4065
rect 13820 4045 13840 4065
rect 13910 4045 13930 4065
rect 14000 4045 14020 4065
rect 14090 4045 14110 4065
rect 14180 4045 14200 4065
rect 14270 4045 14290 4065
rect 14360 4045 14380 4065
rect 14450 4045 14470 4065
rect 14540 4045 14560 4065
rect 14630 4045 14650 4065
rect 14720 4045 14740 4065
rect 14810 4045 14830 4065
rect 14900 4045 14920 4065
rect 14990 4045 15010 4065
rect 15080 4045 15100 4065
rect 15170 4045 15190 4065
rect 15260 4045 15280 4065
rect 15350 4045 15370 4065
rect 15440 4045 15460 4065
rect 15530 4045 15550 4065
rect 15620 4045 15640 4065
rect 15710 4045 15730 4065
rect 15800 4045 15820 4065
rect 15890 4045 15910 4065
rect 15980 4045 16000 4065
rect 16070 4045 16090 4065
rect 16160 4045 16180 4065
rect 16250 4045 16270 4065
rect 16340 4045 16360 4065
rect 16430 4045 16450 4065
rect 16520 4045 16540 4065
rect 16610 4045 16630 4065
rect 16700 4045 16720 4065
rect 16790 4045 16810 4065
rect 16880 4045 16900 4065
rect 16970 4045 16990 4065
rect 17060 4045 17080 4065
rect 17150 4045 17170 4065
rect 17240 4045 17260 4065
rect 17330 4045 17350 4065
rect 17420 4045 17440 4065
rect 17510 4045 17530 4065
rect 17600 4045 17620 4065
rect 17690 4045 17710 4065
rect 17780 4045 17800 4065
rect 17870 4045 17890 4065
rect 17960 4045 17980 4065
rect 18050 4045 18070 4065
rect 18140 4045 18160 4065
rect 18230 4045 18250 4065
rect 18320 4045 18340 4065
rect 18410 4045 18430 4065
rect 18500 4045 18520 4065
rect 18590 4045 18610 4065
rect 18680 4045 18700 4065
rect 18770 4045 18790 4065
rect 18860 4045 18880 4065
rect 18950 4045 18970 4065
rect 19040 4045 19060 4065
rect 19130 4045 19150 4065
rect 19220 4045 19240 4065
rect 19310 4045 19330 4065
rect 19400 4045 19420 4065
rect 19490 4045 19510 4065
rect 19580 4045 19600 4065
rect 19670 4045 19690 4065
rect 19760 4045 19780 4065
rect 19850 4045 19870 4065
rect 19940 4045 19960 4065
rect 20030 4045 20050 4065
rect 20120 4045 20140 4065
rect 20210 4045 20230 4065
rect 20300 4045 20320 4065
rect 20390 4045 20410 4065
rect 20480 4045 20500 4065
rect 20570 4045 20590 4065
rect 20660 4045 20680 4065
rect 9230 3645 9250 3665
rect 9320 3645 9340 3665
rect 9410 3645 9430 3665
rect 9500 3645 9520 3665
rect 9590 3645 9610 3665
rect 9680 3645 9700 3665
rect 9770 3645 9790 3665
rect 9860 3645 9880 3665
rect 9950 3645 9970 3665
rect 10040 3645 10060 3665
rect 10130 3645 10150 3665
rect 10220 3645 10240 3665
rect 10310 3645 10330 3665
rect 10400 3645 10420 3665
rect 10490 3645 10510 3665
rect 10580 3645 10600 3665
rect 10670 3645 10690 3665
rect 10760 3645 10780 3665
rect 10850 3645 10870 3665
rect 10940 3645 10960 3665
rect 11030 3645 11050 3665
rect 11120 3645 11140 3665
rect 11210 3645 11230 3665
rect 11300 3645 11320 3665
rect 11390 3645 11410 3665
rect 11480 3645 11500 3665
rect 11570 3645 11590 3665
rect 11660 3645 11680 3665
rect 11750 3645 11770 3665
rect 11840 3645 11860 3665
rect 11930 3645 11950 3665
rect 12020 3645 12040 3665
rect 12110 3645 12130 3665
rect 12200 3645 12220 3665
rect 12290 3645 12310 3665
rect 12380 3645 12400 3665
rect 12470 3645 12490 3665
rect 12560 3645 12580 3665
rect 12650 3645 12670 3665
rect 12740 3645 12760 3665
rect 12830 3645 12850 3665
rect 12920 3645 12940 3665
rect 13010 3645 13030 3665
rect 13100 3645 13120 3665
rect 13190 3645 13210 3665
rect 13280 3645 13300 3665
rect 13370 3645 13390 3665
rect 13460 3645 13480 3665
rect 13550 3645 13570 3665
rect 13640 3645 13660 3665
rect 13730 3645 13750 3665
rect 13820 3645 13840 3665
rect 13910 3645 13930 3665
rect 14000 3645 14020 3665
rect 14090 3645 14110 3665
rect 14180 3645 14200 3665
rect 14270 3645 14290 3665
rect 14360 3645 14380 3665
rect 14450 3645 14470 3665
rect 14540 3645 14560 3665
rect 14630 3645 14650 3665
rect 14720 3645 14740 3665
rect 14810 3645 14830 3665
rect 14900 3645 14920 3665
rect 14990 3645 15010 3665
rect 15080 3645 15100 3665
rect 15170 3645 15190 3665
rect 15260 3645 15280 3665
rect 15350 3645 15370 3665
rect 15440 3645 15460 3665
rect 15530 3645 15550 3665
rect 15620 3645 15640 3665
rect 15710 3645 15730 3665
rect 15800 3645 15820 3665
rect 15890 3645 15910 3665
rect 15980 3645 16000 3665
rect 16070 3645 16090 3665
rect 16160 3645 16180 3665
rect 16250 3645 16270 3665
rect 16340 3645 16360 3665
rect 16430 3645 16450 3665
rect 16520 3645 16540 3665
rect 16610 3645 16630 3665
rect 16700 3645 16720 3665
rect 16790 3645 16810 3665
rect 16880 3645 16900 3665
rect 16970 3645 16990 3665
rect 17060 3645 17080 3665
rect 17150 3645 17170 3665
rect 17240 3645 17260 3665
rect 17330 3645 17350 3665
rect 17420 3645 17440 3665
rect 17510 3645 17530 3665
rect 17600 3645 17620 3665
rect 17690 3645 17710 3665
rect 17780 3645 17800 3665
rect 17870 3645 17890 3665
rect 17960 3645 17980 3665
rect 18050 3645 18070 3665
rect 18140 3645 18160 3665
rect 18230 3645 18250 3665
rect 18320 3645 18340 3665
rect 18410 3645 18430 3665
rect 18500 3645 18520 3665
rect 18590 3645 18610 3665
rect 18680 3645 18700 3665
rect 18770 3645 18790 3665
rect 18860 3645 18880 3665
rect 18950 3645 18970 3665
rect 19040 3645 19060 3665
rect 19130 3645 19150 3665
rect 19220 3645 19240 3665
rect 19310 3645 19330 3665
rect 19400 3645 19420 3665
rect 19490 3645 19510 3665
rect 19580 3645 19600 3665
rect 19670 3645 19690 3665
rect 19760 3645 19780 3665
rect 19850 3645 19870 3665
rect 19940 3645 19960 3665
rect 20030 3645 20050 3665
rect 20120 3645 20140 3665
rect 20210 3645 20230 3665
rect 20300 3645 20320 3665
rect 20390 3645 20410 3665
rect 20480 3645 20500 3665
rect 20570 3645 20590 3665
rect 20660 3645 20680 3665
rect 9230 3425 9250 3445
rect 9320 3425 9340 3445
rect 9410 3425 9430 3445
rect 9500 3425 9520 3445
rect 9590 3425 9610 3445
rect 9680 3425 9700 3445
rect 9770 3425 9790 3445
rect 9860 3425 9880 3445
rect 9950 3425 9970 3445
rect 10040 3425 10060 3445
rect 10130 3425 10150 3445
rect 10220 3425 10240 3445
rect 10310 3425 10330 3445
rect 10400 3425 10420 3445
rect 10490 3425 10510 3445
rect 10580 3425 10600 3445
rect 10670 3425 10690 3445
rect 10760 3425 10780 3445
rect 10850 3425 10870 3445
rect 10940 3425 10960 3445
rect 11030 3425 11050 3445
rect 11120 3425 11140 3445
rect 11210 3425 11230 3445
rect 11300 3425 11320 3445
rect 11390 3425 11410 3445
rect 11480 3425 11500 3445
rect 11570 3425 11590 3445
rect 11660 3425 11680 3445
rect 11750 3425 11770 3445
rect 11840 3425 11860 3445
rect 11930 3425 11950 3445
rect 12020 3425 12040 3445
rect 12110 3425 12130 3445
rect 12200 3425 12220 3445
rect 12290 3425 12310 3445
rect 12380 3425 12400 3445
rect 12470 3425 12490 3445
rect 12560 3425 12580 3445
rect 12650 3425 12670 3445
rect 12740 3425 12760 3445
rect 12830 3425 12850 3445
rect 12920 3425 12940 3445
rect 13010 3425 13030 3445
rect 13100 3425 13120 3445
rect 13190 3425 13210 3445
rect 13280 3425 13300 3445
rect 13370 3425 13390 3445
rect 13460 3425 13480 3445
rect 13550 3425 13570 3445
rect 13640 3425 13660 3445
rect 13730 3425 13750 3445
rect 13820 3425 13840 3445
rect 13910 3425 13930 3445
rect 14000 3425 14020 3445
rect 14090 3425 14110 3445
rect 14180 3425 14200 3445
rect 14270 3425 14290 3445
rect 14360 3425 14380 3445
rect 14450 3425 14470 3445
rect 14540 3425 14560 3445
rect 14630 3425 14650 3445
rect 14720 3425 14740 3445
rect 14810 3425 14830 3445
rect 14900 3425 14920 3445
rect 14990 3425 15010 3445
rect 15080 3425 15100 3445
rect 15170 3425 15190 3445
rect 15260 3425 15280 3445
rect 15350 3425 15370 3445
rect 15440 3425 15460 3445
rect 15530 3425 15550 3445
rect 15620 3425 15640 3445
rect 15710 3425 15730 3445
rect 15800 3425 15820 3445
rect 15890 3425 15910 3445
rect 15980 3425 16000 3445
rect 16070 3425 16090 3445
rect 16160 3425 16180 3445
rect 16250 3425 16270 3445
rect 16340 3425 16360 3445
rect 16430 3425 16450 3445
rect 16520 3425 16540 3445
rect 16610 3425 16630 3445
rect 16700 3425 16720 3445
rect 16790 3425 16810 3445
rect 16880 3425 16900 3445
rect 16970 3425 16990 3445
rect 17060 3425 17080 3445
rect 17150 3425 17170 3445
rect 17240 3425 17260 3445
rect 17330 3425 17350 3445
rect 17420 3425 17440 3445
rect 17510 3425 17530 3445
rect 17600 3425 17620 3445
rect 17690 3425 17710 3445
rect 17780 3425 17800 3445
rect 17870 3425 17890 3445
rect 17960 3425 17980 3445
rect 18050 3425 18070 3445
rect 18140 3425 18160 3445
rect 18230 3425 18250 3445
rect 18320 3425 18340 3445
rect 18410 3425 18430 3445
rect 18500 3425 18520 3445
rect 18590 3425 18610 3445
rect 18680 3425 18700 3445
rect 18770 3425 18790 3445
rect 18860 3425 18880 3445
rect 18950 3425 18970 3445
rect 19040 3425 19060 3445
rect 19130 3425 19150 3445
rect 19220 3425 19240 3445
rect 19310 3425 19330 3445
rect 19400 3425 19420 3445
rect 19490 3425 19510 3445
rect 19580 3425 19600 3445
rect 19670 3425 19690 3445
rect 19760 3425 19780 3445
rect 19850 3425 19870 3445
rect 19940 3425 19960 3445
rect 20030 3425 20050 3445
rect 20120 3425 20140 3445
rect 20210 3425 20230 3445
rect 20300 3425 20320 3445
rect 20390 3425 20410 3445
rect 20480 3425 20500 3445
rect 20570 3425 20590 3445
rect 20660 3425 20680 3445
<< nsubdiffcont >>
rect 9230 4345 9250 4365
rect 9320 4345 9340 4365
rect 9410 4345 9430 4365
rect 9500 4345 9520 4365
rect 9590 4345 9610 4365
rect 9680 4345 9700 4365
rect 9770 4345 9790 4365
rect 9860 4345 9880 4365
rect 9950 4345 9970 4365
rect 10040 4345 10060 4365
rect 10130 4345 10150 4365
rect 10220 4345 10240 4365
rect 10310 4345 10330 4365
rect 10400 4345 10420 4365
rect 10490 4345 10510 4365
rect 10580 4345 10600 4365
rect 10670 4345 10690 4365
rect 10760 4345 10780 4365
rect 10850 4345 10870 4365
rect 10940 4345 10960 4365
rect 11030 4345 11050 4365
rect 11120 4345 11140 4365
rect 11210 4345 11230 4365
rect 11300 4345 11320 4365
rect 11390 4345 11410 4365
rect 11480 4345 11500 4365
rect 11570 4345 11590 4365
rect 11660 4345 11680 4365
rect 11750 4345 11770 4365
rect 11840 4345 11860 4365
rect 11930 4345 11950 4365
rect 12020 4345 12040 4365
rect 12110 4345 12130 4365
rect 12200 4345 12220 4365
rect 12290 4345 12310 4365
rect 12380 4345 12400 4365
rect 12470 4345 12490 4365
rect 12560 4345 12580 4365
rect 12650 4345 12670 4365
rect 12740 4345 12760 4365
rect 12830 4345 12850 4365
rect 12920 4345 12940 4365
rect 13010 4345 13030 4365
rect 13100 4345 13120 4365
rect 13190 4345 13210 4365
rect 13280 4345 13300 4365
rect 13370 4345 13390 4365
rect 13460 4345 13480 4365
rect 13550 4345 13570 4365
rect 13640 4345 13660 4365
rect 13730 4345 13750 4365
rect 13820 4345 13840 4365
rect 13910 4345 13930 4365
rect 14000 4345 14020 4365
rect 14090 4345 14110 4365
rect 14180 4345 14200 4365
rect 14270 4345 14290 4365
rect 14360 4345 14380 4365
rect 14450 4345 14470 4365
rect 14540 4345 14560 4365
rect 14630 4345 14650 4365
rect 14720 4345 14740 4365
rect 14810 4345 14830 4365
rect 14900 4345 14920 4365
rect 14990 4345 15010 4365
rect 15080 4345 15100 4365
rect 15170 4345 15190 4365
rect 15260 4345 15280 4365
rect 15350 4345 15370 4365
rect 15440 4345 15460 4365
rect 15530 4345 15550 4365
rect 15620 4345 15640 4365
rect 15710 4345 15730 4365
rect 15800 4345 15820 4365
rect 15890 4345 15910 4365
rect 15980 4345 16000 4365
rect 16070 4345 16090 4365
rect 16160 4345 16180 4365
rect 16250 4345 16270 4365
rect 16340 4345 16360 4365
rect 16430 4345 16450 4365
rect 16520 4345 16540 4365
rect 16610 4345 16630 4365
rect 16700 4345 16720 4365
rect 16790 4345 16810 4365
rect 16880 4345 16900 4365
rect 16970 4345 16990 4365
rect 17060 4345 17080 4365
rect 17150 4345 17170 4365
rect 17240 4345 17260 4365
rect 17330 4345 17350 4365
rect 17420 4345 17440 4365
rect 17510 4345 17530 4365
rect 17600 4345 17620 4365
rect 17690 4345 17710 4365
rect 17780 4345 17800 4365
rect 17870 4345 17890 4365
rect 17960 4345 17980 4365
rect 18050 4345 18070 4365
rect 18140 4345 18160 4365
rect 18230 4345 18250 4365
rect 18320 4345 18340 4365
rect 18410 4345 18430 4365
rect 18500 4345 18520 4365
rect 18590 4345 18610 4365
rect 18680 4345 18700 4365
rect 18770 4345 18790 4365
rect 18860 4345 18880 4365
rect 18950 4345 18970 4365
rect 19040 4345 19060 4365
rect 19130 4345 19150 4365
rect 19220 4345 19240 4365
rect 19310 4345 19330 4365
rect 19400 4345 19420 4365
rect 19490 4345 19510 4365
rect 19580 4345 19600 4365
rect 19670 4345 19690 4365
rect 19760 4345 19780 4365
rect 19850 4345 19870 4365
rect 19940 4345 19960 4365
rect 20030 4345 20050 4365
rect 20120 4345 20140 4365
rect 20210 4345 20230 4365
rect 20300 4345 20320 4365
rect 20390 4345 20410 4365
rect 20480 4345 20500 4365
rect 20570 4345 20590 4365
rect 20660 4345 20680 4365
rect 9230 4125 9250 4145
rect 9320 4125 9340 4145
rect 9410 4125 9430 4145
rect 9500 4125 9520 4145
rect 9590 4125 9610 4145
rect 9680 4125 9700 4145
rect 9770 4125 9790 4145
rect 9860 4125 9880 4145
rect 9950 4125 9970 4145
rect 10040 4125 10060 4145
rect 10130 4125 10150 4145
rect 10220 4125 10240 4145
rect 10310 4125 10330 4145
rect 10400 4125 10420 4145
rect 10490 4125 10510 4145
rect 10580 4125 10600 4145
rect 10670 4125 10690 4145
rect 10760 4125 10780 4145
rect 10850 4125 10870 4145
rect 10940 4125 10960 4145
rect 11030 4125 11050 4145
rect 11120 4125 11140 4145
rect 11210 4125 11230 4145
rect 11300 4125 11320 4145
rect 11390 4125 11410 4145
rect 11480 4125 11500 4145
rect 11570 4125 11590 4145
rect 11660 4125 11680 4145
rect 11750 4125 11770 4145
rect 11840 4125 11860 4145
rect 11930 4125 11950 4145
rect 12020 4125 12040 4145
rect 12110 4125 12130 4145
rect 12200 4125 12220 4145
rect 12290 4125 12310 4145
rect 12380 4125 12400 4145
rect 12470 4125 12490 4145
rect 12560 4125 12580 4145
rect 12650 4125 12670 4145
rect 12740 4125 12760 4145
rect 12830 4125 12850 4145
rect 12920 4125 12940 4145
rect 13010 4125 13030 4145
rect 13100 4125 13120 4145
rect 13190 4125 13210 4145
rect 13280 4125 13300 4145
rect 13370 4125 13390 4145
rect 13460 4125 13480 4145
rect 13550 4125 13570 4145
rect 13640 4125 13660 4145
rect 13730 4125 13750 4145
rect 13820 4125 13840 4145
rect 13910 4125 13930 4145
rect 14000 4125 14020 4145
rect 14090 4125 14110 4145
rect 14180 4125 14200 4145
rect 14270 4125 14290 4145
rect 14360 4125 14380 4145
rect 14450 4125 14470 4145
rect 14540 4125 14560 4145
rect 14630 4125 14650 4145
rect 14720 4125 14740 4145
rect 14810 4125 14830 4145
rect 14900 4125 14920 4145
rect 14990 4125 15010 4145
rect 15080 4125 15100 4145
rect 15170 4125 15190 4145
rect 15260 4125 15280 4145
rect 15350 4125 15370 4145
rect 15440 4125 15460 4145
rect 15530 4125 15550 4145
rect 15620 4125 15640 4145
rect 15710 4125 15730 4145
rect 15800 4125 15820 4145
rect 15890 4125 15910 4145
rect 15980 4125 16000 4145
rect 16070 4125 16090 4145
rect 16160 4125 16180 4145
rect 16250 4125 16270 4145
rect 16340 4125 16360 4145
rect 16430 4125 16450 4145
rect 16520 4125 16540 4145
rect 16610 4125 16630 4145
rect 16700 4125 16720 4145
rect 16790 4125 16810 4145
rect 16880 4125 16900 4145
rect 16970 4125 16990 4145
rect 17060 4125 17080 4145
rect 17150 4125 17170 4145
rect 17240 4125 17260 4145
rect 17330 4125 17350 4145
rect 17420 4125 17440 4145
rect 17510 4125 17530 4145
rect 17600 4125 17620 4145
rect 17690 4125 17710 4145
rect 17780 4125 17800 4145
rect 17870 4125 17890 4145
rect 17960 4125 17980 4145
rect 18050 4125 18070 4145
rect 18140 4125 18160 4145
rect 18230 4125 18250 4145
rect 18320 4125 18340 4145
rect 18410 4125 18430 4145
rect 18500 4125 18520 4145
rect 18590 4125 18610 4145
rect 18680 4125 18700 4145
rect 18770 4125 18790 4145
rect 18860 4125 18880 4145
rect 18950 4125 18970 4145
rect 19040 4125 19060 4145
rect 19130 4125 19150 4145
rect 19220 4125 19240 4145
rect 19310 4125 19330 4145
rect 19400 4125 19420 4145
rect 19490 4125 19510 4145
rect 19580 4125 19600 4145
rect 19670 4125 19690 4145
rect 19760 4125 19780 4145
rect 19850 4125 19870 4145
rect 19940 4125 19960 4145
rect 20030 4125 20050 4145
rect 20120 4125 20140 4145
rect 20210 4125 20230 4145
rect 20300 4125 20320 4145
rect 20390 4125 20410 4145
rect 20480 4125 20500 4145
rect 20570 4125 20590 4145
rect 20660 4125 20680 4145
<< poly >>
rect 9215 4315 9265 4330
rect 9305 4315 9355 4330
rect 9395 4315 9445 4330
rect 9485 4315 9535 4330
rect 9575 4315 9625 4330
rect 9665 4315 9715 4330
rect 9755 4315 9805 4330
rect 9845 4315 9895 4330
rect 9935 4315 9985 4330
rect 10025 4315 10075 4330
rect 10115 4315 10165 4330
rect 10205 4315 10255 4330
rect 10295 4315 10345 4330
rect 10385 4315 10435 4330
rect 10475 4315 10525 4330
rect 10565 4315 10615 4330
rect 10655 4315 10705 4330
rect 10745 4315 10795 4330
rect 10835 4315 10885 4330
rect 10925 4315 10975 4330
rect 11015 4315 11065 4330
rect 11105 4315 11155 4330
rect 11195 4315 11245 4330
rect 11285 4315 11335 4330
rect 11375 4315 11425 4330
rect 11465 4315 11515 4330
rect 11555 4315 11605 4330
rect 11645 4315 11695 4330
rect 11735 4315 11785 4330
rect 11825 4315 11875 4330
rect 11915 4315 11965 4330
rect 12005 4315 12055 4330
rect 12095 4315 12145 4330
rect 12185 4315 12235 4330
rect 12275 4315 12325 4330
rect 12365 4315 12415 4330
rect 12455 4315 12505 4330
rect 12545 4315 12595 4330
rect 12635 4315 12685 4330
rect 12725 4315 12775 4330
rect 12815 4315 12865 4330
rect 12905 4315 12955 4330
rect 12995 4315 13045 4330
rect 13085 4315 13135 4330
rect 13175 4315 13225 4330
rect 13265 4315 13315 4330
rect 13355 4315 13405 4330
rect 13445 4315 13495 4330
rect 13535 4315 13585 4330
rect 13625 4315 13675 4330
rect 13715 4315 13765 4330
rect 13805 4315 13855 4330
rect 13895 4315 13945 4330
rect 13985 4315 14035 4330
rect 14075 4315 14125 4330
rect 14165 4315 14215 4330
rect 14255 4315 14305 4330
rect 14345 4315 14395 4330
rect 14435 4315 14485 4330
rect 14525 4315 14575 4330
rect 14615 4315 14665 4330
rect 14705 4315 14755 4330
rect 14795 4315 14845 4330
rect 14885 4315 14935 4330
rect 14975 4315 15025 4330
rect 15065 4315 15115 4330
rect 15155 4315 15205 4330
rect 15245 4315 15295 4330
rect 15335 4315 15385 4330
rect 15425 4315 15475 4330
rect 15515 4315 15565 4330
rect 15605 4315 15655 4330
rect 15695 4315 15745 4330
rect 15785 4315 15835 4330
rect 15875 4315 15925 4330
rect 15965 4315 16015 4330
rect 16055 4315 16105 4330
rect 16145 4315 16195 4330
rect 16235 4315 16285 4330
rect 16325 4315 16375 4330
rect 16415 4315 16465 4330
rect 16505 4315 16555 4330
rect 16595 4315 16645 4330
rect 16685 4315 16735 4330
rect 16775 4315 16825 4330
rect 16865 4315 16915 4330
rect 16955 4315 17005 4330
rect 17045 4315 17095 4330
rect 17135 4315 17185 4330
rect 17225 4315 17275 4330
rect 17315 4315 17365 4330
rect 17405 4315 17455 4330
rect 17495 4315 17545 4330
rect 17585 4315 17635 4330
rect 17675 4315 17725 4330
rect 17765 4315 17815 4330
rect 17855 4315 17905 4330
rect 17945 4315 17995 4330
rect 18035 4315 18085 4330
rect 18125 4315 18175 4330
rect 18215 4315 18265 4330
rect 18305 4315 18355 4330
rect 18395 4315 18445 4330
rect 18485 4315 18535 4330
rect 18575 4315 18625 4330
rect 18665 4315 18715 4330
rect 18755 4315 18805 4330
rect 18845 4315 18895 4330
rect 18935 4315 18985 4330
rect 19025 4315 19075 4330
rect 19115 4315 19165 4330
rect 19205 4315 19255 4330
rect 19295 4315 19345 4330
rect 19385 4315 19435 4330
rect 19475 4315 19525 4330
rect 19565 4315 19615 4330
rect 19655 4315 19705 4330
rect 19745 4315 19795 4330
rect 19835 4315 19885 4330
rect 19925 4315 19975 4330
rect 20015 4315 20065 4330
rect 20105 4315 20155 4330
rect 20195 4315 20245 4330
rect 20285 4315 20335 4330
rect 20375 4315 20425 4330
rect 20465 4315 20515 4330
rect 20555 4315 20605 4330
rect 20645 4315 20695 4330
rect 9215 4195 9265 4215
rect 9305 4195 9355 4215
rect 9215 4190 9355 4195
rect 9215 4170 9230 4190
rect 9250 4170 9320 4190
rect 9340 4170 9355 4190
rect 9215 4165 9355 4170
rect 9395 4195 9445 4215
rect 9485 4195 9535 4215
rect 9395 4190 9535 4195
rect 9395 4170 9410 4190
rect 9430 4170 9500 4190
rect 9520 4170 9535 4190
rect 9395 4165 9535 4170
rect 9575 4195 9625 4215
rect 9665 4195 9715 4215
rect 9575 4190 9715 4195
rect 9575 4170 9590 4190
rect 9610 4170 9680 4190
rect 9700 4170 9715 4190
rect 9575 4165 9715 4170
rect 9755 4195 9805 4215
rect 9845 4195 9895 4215
rect 9755 4190 9895 4195
rect 9755 4170 9770 4190
rect 9790 4170 9860 4190
rect 9880 4170 9895 4190
rect 9755 4165 9895 4170
rect 9935 4195 9985 4215
rect 10025 4195 10075 4215
rect 9935 4190 10075 4195
rect 9935 4170 9950 4190
rect 9970 4170 10040 4190
rect 10060 4170 10075 4190
rect 9935 4165 10075 4170
rect 10115 4195 10165 4215
rect 10205 4195 10255 4215
rect 10115 4190 10255 4195
rect 10115 4170 10130 4190
rect 10150 4170 10220 4190
rect 10240 4170 10255 4190
rect 10115 4165 10255 4170
rect 10295 4195 10345 4215
rect 10385 4195 10435 4215
rect 10295 4190 10435 4195
rect 10295 4170 10310 4190
rect 10330 4170 10400 4190
rect 10420 4170 10435 4190
rect 10295 4165 10435 4170
rect 10475 4195 10525 4215
rect 10565 4195 10615 4215
rect 10475 4190 10615 4195
rect 10475 4170 10490 4190
rect 10510 4170 10580 4190
rect 10600 4170 10615 4190
rect 10475 4165 10615 4170
rect 10655 4195 10705 4215
rect 10745 4195 10795 4215
rect 10655 4190 10795 4195
rect 10655 4170 10670 4190
rect 10690 4170 10760 4190
rect 10780 4170 10795 4190
rect 10655 4165 10795 4170
rect 10835 4195 10885 4215
rect 10925 4195 10975 4215
rect 10835 4190 10975 4195
rect 10835 4170 10850 4190
rect 10870 4170 10940 4190
rect 10960 4170 10975 4190
rect 10835 4165 10975 4170
rect 11015 4195 11065 4215
rect 11105 4195 11155 4215
rect 11015 4190 11155 4195
rect 11015 4170 11030 4190
rect 11050 4170 11120 4190
rect 11140 4170 11155 4190
rect 11015 4165 11155 4170
rect 11195 4195 11245 4215
rect 11285 4195 11335 4215
rect 11195 4190 11335 4195
rect 11195 4170 11210 4190
rect 11230 4170 11300 4190
rect 11320 4170 11335 4190
rect 11195 4165 11335 4170
rect 11375 4195 11425 4215
rect 11465 4195 11515 4215
rect 11375 4190 11515 4195
rect 11375 4170 11390 4190
rect 11410 4170 11480 4190
rect 11500 4170 11515 4190
rect 11375 4165 11515 4170
rect 11555 4195 11605 4215
rect 11645 4195 11695 4215
rect 11555 4190 11695 4195
rect 11555 4170 11570 4190
rect 11590 4170 11660 4190
rect 11680 4170 11695 4190
rect 11555 4165 11695 4170
rect 11735 4195 11785 4215
rect 11825 4195 11875 4215
rect 11735 4190 11875 4195
rect 11735 4170 11750 4190
rect 11770 4170 11840 4190
rect 11860 4170 11875 4190
rect 11735 4165 11875 4170
rect 11915 4195 11965 4215
rect 12005 4195 12055 4215
rect 11915 4190 12055 4195
rect 11915 4170 11930 4190
rect 11950 4170 12020 4190
rect 12040 4170 12055 4190
rect 11915 4165 12055 4170
rect 12095 4195 12145 4215
rect 12185 4195 12235 4215
rect 12095 4190 12235 4195
rect 12095 4170 12110 4190
rect 12130 4170 12200 4190
rect 12220 4170 12235 4190
rect 12095 4165 12235 4170
rect 12275 4195 12325 4215
rect 12365 4195 12415 4215
rect 12275 4190 12415 4195
rect 12275 4170 12290 4190
rect 12310 4170 12380 4190
rect 12400 4170 12415 4190
rect 12275 4165 12415 4170
rect 12455 4195 12505 4215
rect 12545 4195 12595 4215
rect 12455 4190 12595 4195
rect 12455 4170 12470 4190
rect 12490 4170 12560 4190
rect 12580 4170 12595 4190
rect 12455 4165 12595 4170
rect 12635 4195 12685 4215
rect 12725 4195 12775 4215
rect 12635 4190 12775 4195
rect 12635 4170 12650 4190
rect 12670 4170 12740 4190
rect 12760 4170 12775 4190
rect 12635 4165 12775 4170
rect 12815 4195 12865 4215
rect 12905 4195 12955 4215
rect 12815 4190 12955 4195
rect 12815 4170 12830 4190
rect 12850 4170 12920 4190
rect 12940 4170 12955 4190
rect 12815 4165 12955 4170
rect 12995 4195 13045 4215
rect 13085 4195 13135 4215
rect 12995 4190 13135 4195
rect 12995 4170 13010 4190
rect 13030 4170 13100 4190
rect 13120 4170 13135 4190
rect 12995 4165 13135 4170
rect 13175 4195 13225 4215
rect 13265 4195 13315 4215
rect 13175 4190 13315 4195
rect 13175 4170 13190 4190
rect 13210 4170 13280 4190
rect 13300 4170 13315 4190
rect 13175 4165 13315 4170
rect 13355 4195 13405 4215
rect 13445 4195 13495 4215
rect 13355 4190 13495 4195
rect 13355 4170 13370 4190
rect 13390 4170 13460 4190
rect 13480 4170 13495 4190
rect 13355 4165 13495 4170
rect 13535 4195 13585 4215
rect 13625 4195 13675 4215
rect 13535 4190 13675 4195
rect 13535 4170 13550 4190
rect 13570 4170 13640 4190
rect 13660 4170 13675 4190
rect 13535 4165 13675 4170
rect 13715 4195 13765 4215
rect 13805 4195 13855 4215
rect 13715 4190 13855 4195
rect 13715 4170 13730 4190
rect 13750 4170 13820 4190
rect 13840 4170 13855 4190
rect 13715 4165 13855 4170
rect 13895 4195 13945 4215
rect 13985 4195 14035 4215
rect 13895 4190 14035 4195
rect 13895 4170 13910 4190
rect 13930 4170 14000 4190
rect 14020 4170 14035 4190
rect 13895 4165 14035 4170
rect 14075 4195 14125 4215
rect 14165 4195 14215 4215
rect 14075 4190 14215 4195
rect 14075 4170 14090 4190
rect 14110 4170 14180 4190
rect 14200 4170 14215 4190
rect 14075 4165 14215 4170
rect 14255 4195 14305 4215
rect 14345 4195 14395 4215
rect 14255 4190 14395 4195
rect 14255 4170 14270 4190
rect 14290 4170 14360 4190
rect 14380 4170 14395 4190
rect 14255 4165 14395 4170
rect 14435 4195 14485 4215
rect 14525 4195 14575 4215
rect 14435 4190 14575 4195
rect 14435 4170 14450 4190
rect 14470 4170 14540 4190
rect 14560 4170 14575 4190
rect 14435 4165 14575 4170
rect 14615 4195 14665 4215
rect 14705 4195 14755 4215
rect 14615 4190 14755 4195
rect 14615 4170 14630 4190
rect 14650 4170 14720 4190
rect 14740 4170 14755 4190
rect 14615 4165 14755 4170
rect 14795 4195 14845 4215
rect 14885 4195 14935 4215
rect 14795 4190 14935 4195
rect 14795 4170 14810 4190
rect 14830 4170 14900 4190
rect 14920 4170 14935 4190
rect 14795 4165 14935 4170
rect 14975 4195 15025 4215
rect 15065 4195 15115 4215
rect 14975 4190 15115 4195
rect 14975 4170 14990 4190
rect 15010 4170 15080 4190
rect 15100 4170 15115 4190
rect 14975 4165 15115 4170
rect 15155 4195 15205 4215
rect 15245 4195 15295 4215
rect 15155 4190 15295 4195
rect 15155 4170 15170 4190
rect 15190 4170 15260 4190
rect 15280 4170 15295 4190
rect 15155 4165 15295 4170
rect 15335 4195 15385 4215
rect 15425 4195 15475 4215
rect 15335 4190 15475 4195
rect 15335 4170 15350 4190
rect 15370 4170 15440 4190
rect 15460 4170 15475 4190
rect 15335 4165 15475 4170
rect 15515 4195 15565 4215
rect 15605 4195 15655 4215
rect 15515 4190 15655 4195
rect 15515 4170 15530 4190
rect 15550 4170 15620 4190
rect 15640 4170 15655 4190
rect 15515 4165 15655 4170
rect 15695 4195 15745 4215
rect 15785 4195 15835 4215
rect 15695 4190 15835 4195
rect 15695 4170 15710 4190
rect 15730 4170 15800 4190
rect 15820 4170 15835 4190
rect 15695 4165 15835 4170
rect 15875 4195 15925 4215
rect 15965 4195 16015 4215
rect 15875 4190 16015 4195
rect 15875 4170 15890 4190
rect 15910 4170 15980 4190
rect 16000 4170 16015 4190
rect 15875 4165 16015 4170
rect 16055 4195 16105 4215
rect 16145 4195 16195 4215
rect 16055 4190 16195 4195
rect 16055 4170 16070 4190
rect 16090 4170 16160 4190
rect 16180 4170 16195 4190
rect 16055 4165 16195 4170
rect 16235 4195 16285 4215
rect 16325 4195 16375 4215
rect 16235 4190 16375 4195
rect 16235 4170 16250 4190
rect 16270 4170 16340 4190
rect 16360 4170 16375 4190
rect 16235 4165 16375 4170
rect 16415 4195 16465 4215
rect 16505 4195 16555 4215
rect 16415 4190 16555 4195
rect 16415 4170 16430 4190
rect 16450 4170 16520 4190
rect 16540 4170 16555 4190
rect 16415 4165 16555 4170
rect 16595 4195 16645 4215
rect 16685 4195 16735 4215
rect 16595 4190 16735 4195
rect 16595 4170 16610 4190
rect 16630 4170 16700 4190
rect 16720 4170 16735 4190
rect 16595 4165 16735 4170
rect 16775 4195 16825 4215
rect 16865 4195 16915 4215
rect 16775 4190 16915 4195
rect 16775 4170 16790 4190
rect 16810 4170 16880 4190
rect 16900 4170 16915 4190
rect 16775 4165 16915 4170
rect 16955 4195 17005 4215
rect 17045 4195 17095 4215
rect 16955 4190 17095 4195
rect 16955 4170 16970 4190
rect 16990 4170 17060 4190
rect 17080 4170 17095 4190
rect 16955 4165 17095 4170
rect 17135 4195 17185 4215
rect 17225 4195 17275 4215
rect 17135 4190 17275 4195
rect 17135 4170 17150 4190
rect 17170 4170 17240 4190
rect 17260 4170 17275 4190
rect 17135 4165 17275 4170
rect 17315 4195 17365 4215
rect 17405 4195 17455 4215
rect 17315 4190 17455 4195
rect 17315 4170 17330 4190
rect 17350 4170 17420 4190
rect 17440 4170 17455 4190
rect 17315 4165 17455 4170
rect 17495 4195 17545 4215
rect 17585 4195 17635 4215
rect 17495 4190 17635 4195
rect 17495 4170 17510 4190
rect 17530 4170 17600 4190
rect 17620 4170 17635 4190
rect 17495 4165 17635 4170
rect 17675 4195 17725 4215
rect 17765 4195 17815 4215
rect 17675 4190 17815 4195
rect 17675 4170 17690 4190
rect 17710 4170 17780 4190
rect 17800 4170 17815 4190
rect 17675 4165 17815 4170
rect 17855 4195 17905 4215
rect 17945 4195 17995 4215
rect 17855 4190 17995 4195
rect 17855 4170 17870 4190
rect 17890 4170 17960 4190
rect 17980 4170 17995 4190
rect 17855 4165 17995 4170
rect 18035 4195 18085 4215
rect 18125 4195 18175 4215
rect 18035 4190 18175 4195
rect 18035 4170 18050 4190
rect 18070 4170 18140 4190
rect 18160 4170 18175 4190
rect 18035 4165 18175 4170
rect 18215 4195 18265 4215
rect 18305 4195 18355 4215
rect 18215 4190 18355 4195
rect 18215 4170 18230 4190
rect 18250 4170 18320 4190
rect 18340 4170 18355 4190
rect 18215 4165 18355 4170
rect 18395 4195 18445 4215
rect 18485 4195 18535 4215
rect 18395 4190 18535 4195
rect 18395 4170 18410 4190
rect 18430 4170 18500 4190
rect 18520 4170 18535 4190
rect 18395 4165 18535 4170
rect 18575 4195 18625 4215
rect 18665 4195 18715 4215
rect 18575 4190 18715 4195
rect 18575 4170 18590 4190
rect 18610 4170 18680 4190
rect 18700 4170 18715 4190
rect 18575 4165 18715 4170
rect 18755 4195 18805 4215
rect 18845 4195 18895 4215
rect 18755 4190 18895 4195
rect 18755 4170 18770 4190
rect 18790 4170 18860 4190
rect 18880 4170 18895 4190
rect 18755 4165 18895 4170
rect 18935 4195 18985 4215
rect 19025 4195 19075 4215
rect 18935 4190 19075 4195
rect 18935 4170 18950 4190
rect 18970 4170 19040 4190
rect 19060 4170 19075 4190
rect 18935 4165 19075 4170
rect 19115 4195 19165 4215
rect 19205 4195 19255 4215
rect 19115 4190 19255 4195
rect 19115 4170 19130 4190
rect 19150 4170 19220 4190
rect 19240 4170 19255 4190
rect 19115 4165 19255 4170
rect 19295 4195 19345 4215
rect 19385 4195 19435 4215
rect 19295 4190 19435 4195
rect 19295 4170 19310 4190
rect 19330 4170 19400 4190
rect 19420 4170 19435 4190
rect 19295 4165 19435 4170
rect 19475 4195 19525 4215
rect 19565 4195 19615 4215
rect 19475 4190 19615 4195
rect 19475 4170 19490 4190
rect 19510 4170 19580 4190
rect 19600 4170 19615 4190
rect 19475 4165 19615 4170
rect 19655 4195 19705 4215
rect 19745 4195 19795 4215
rect 19655 4190 19795 4195
rect 19655 4170 19670 4190
rect 19690 4170 19760 4190
rect 19780 4170 19795 4190
rect 19655 4165 19795 4170
rect 19835 4195 19885 4215
rect 19925 4195 19975 4215
rect 19835 4190 19975 4195
rect 19835 4170 19850 4190
rect 19870 4170 19940 4190
rect 19960 4170 19975 4190
rect 19835 4165 19975 4170
rect 20015 4195 20065 4215
rect 20105 4195 20155 4215
rect 20015 4190 20155 4195
rect 20015 4170 20030 4190
rect 20050 4170 20120 4190
rect 20140 4170 20155 4190
rect 20015 4165 20155 4170
rect 20195 4195 20245 4215
rect 20285 4195 20335 4215
rect 20195 4190 20335 4195
rect 20195 4170 20210 4190
rect 20230 4170 20300 4190
rect 20320 4170 20335 4190
rect 20195 4165 20335 4170
rect 20375 4195 20425 4215
rect 20465 4195 20515 4215
rect 20375 4190 20515 4195
rect 20375 4170 20390 4190
rect 20410 4170 20480 4190
rect 20500 4170 20515 4190
rect 20375 4165 20515 4170
rect 20555 4195 20605 4215
rect 20645 4195 20695 4215
rect 20555 4190 20695 4195
rect 20555 4170 20570 4190
rect 20590 4170 20660 4190
rect 20680 4170 20695 4190
rect 20555 4165 20695 4170
rect 9215 3620 9355 3625
rect 9215 3600 9230 3620
rect 9250 3600 9320 3620
rect 9340 3600 9355 3620
rect 9215 3595 9355 3600
rect 9215 3575 9265 3595
rect 9305 3575 9355 3595
rect 9395 3620 9535 3625
rect 9395 3600 9410 3620
rect 9430 3600 9500 3620
rect 9520 3600 9535 3620
rect 9395 3595 9535 3600
rect 9395 3575 9445 3595
rect 9485 3575 9535 3595
rect 9575 3620 9715 3625
rect 9575 3600 9590 3620
rect 9610 3600 9680 3620
rect 9700 3600 9715 3620
rect 9575 3595 9715 3600
rect 9575 3575 9625 3595
rect 9665 3575 9715 3595
rect 9755 3620 9895 3625
rect 9755 3600 9770 3620
rect 9790 3600 9860 3620
rect 9880 3600 9895 3620
rect 9755 3595 9895 3600
rect 9755 3575 9805 3595
rect 9845 3575 9895 3595
rect 9935 3620 10075 3625
rect 9935 3600 9950 3620
rect 9970 3600 10040 3620
rect 10060 3600 10075 3620
rect 9935 3595 10075 3600
rect 9935 3575 9985 3595
rect 10025 3575 10075 3595
rect 10115 3620 10255 3625
rect 10115 3600 10130 3620
rect 10150 3600 10220 3620
rect 10240 3600 10255 3620
rect 10115 3595 10255 3600
rect 10115 3575 10165 3595
rect 10205 3575 10255 3595
rect 10295 3620 10435 3625
rect 10295 3600 10310 3620
rect 10330 3600 10400 3620
rect 10420 3600 10435 3620
rect 10295 3595 10435 3600
rect 10295 3575 10345 3595
rect 10385 3575 10435 3595
rect 10475 3620 10615 3625
rect 10475 3600 10490 3620
rect 10510 3600 10580 3620
rect 10600 3600 10615 3620
rect 10475 3595 10615 3600
rect 10475 3575 10525 3595
rect 10565 3575 10615 3595
rect 10655 3620 10795 3625
rect 10655 3600 10670 3620
rect 10690 3600 10760 3620
rect 10780 3600 10795 3620
rect 10655 3595 10795 3600
rect 10655 3575 10705 3595
rect 10745 3575 10795 3595
rect 10835 3620 10975 3625
rect 10835 3600 10850 3620
rect 10870 3600 10940 3620
rect 10960 3600 10975 3620
rect 10835 3595 10975 3600
rect 10835 3575 10885 3595
rect 10925 3575 10975 3595
rect 11015 3620 11155 3625
rect 11015 3600 11030 3620
rect 11050 3600 11120 3620
rect 11140 3600 11155 3620
rect 11015 3595 11155 3600
rect 11015 3575 11065 3595
rect 11105 3575 11155 3595
rect 11195 3620 11335 3625
rect 11195 3600 11210 3620
rect 11230 3600 11300 3620
rect 11320 3600 11335 3620
rect 11195 3595 11335 3600
rect 11195 3575 11245 3595
rect 11285 3575 11335 3595
rect 11375 3620 11515 3625
rect 11375 3600 11390 3620
rect 11410 3600 11480 3620
rect 11500 3600 11515 3620
rect 11375 3595 11515 3600
rect 11375 3575 11425 3595
rect 11465 3575 11515 3595
rect 11555 3620 11695 3625
rect 11555 3600 11570 3620
rect 11590 3600 11660 3620
rect 11680 3600 11695 3620
rect 11555 3595 11695 3600
rect 11555 3575 11605 3595
rect 11645 3575 11695 3595
rect 11735 3620 11875 3625
rect 11735 3600 11750 3620
rect 11770 3600 11840 3620
rect 11860 3600 11875 3620
rect 11735 3595 11875 3600
rect 11735 3575 11785 3595
rect 11825 3575 11875 3595
rect 11915 3620 12055 3625
rect 11915 3600 11930 3620
rect 11950 3600 12020 3620
rect 12040 3600 12055 3620
rect 11915 3595 12055 3600
rect 11915 3575 11965 3595
rect 12005 3575 12055 3595
rect 12095 3620 12235 3625
rect 12095 3600 12110 3620
rect 12130 3600 12200 3620
rect 12220 3600 12235 3620
rect 12095 3595 12235 3600
rect 12095 3575 12145 3595
rect 12185 3575 12235 3595
rect 12275 3620 12415 3625
rect 12275 3600 12290 3620
rect 12310 3600 12380 3620
rect 12400 3600 12415 3620
rect 12275 3595 12415 3600
rect 12275 3575 12325 3595
rect 12365 3575 12415 3595
rect 12455 3620 12595 3625
rect 12455 3600 12470 3620
rect 12490 3600 12560 3620
rect 12580 3600 12595 3620
rect 12455 3595 12595 3600
rect 12455 3575 12505 3595
rect 12545 3575 12595 3595
rect 12635 3620 12775 3625
rect 12635 3600 12650 3620
rect 12670 3600 12740 3620
rect 12760 3600 12775 3620
rect 12635 3595 12775 3600
rect 12635 3575 12685 3595
rect 12725 3575 12775 3595
rect 12815 3620 12955 3625
rect 12815 3600 12830 3620
rect 12850 3600 12920 3620
rect 12940 3600 12955 3620
rect 12815 3595 12955 3600
rect 12815 3575 12865 3595
rect 12905 3575 12955 3595
rect 12995 3620 13135 3625
rect 12995 3600 13010 3620
rect 13030 3600 13100 3620
rect 13120 3600 13135 3620
rect 12995 3595 13135 3600
rect 12995 3575 13045 3595
rect 13085 3575 13135 3595
rect 13175 3620 13315 3625
rect 13175 3600 13190 3620
rect 13210 3600 13280 3620
rect 13300 3600 13315 3620
rect 13175 3595 13315 3600
rect 13175 3575 13225 3595
rect 13265 3575 13315 3595
rect 13355 3620 13495 3625
rect 13355 3600 13370 3620
rect 13390 3600 13460 3620
rect 13480 3600 13495 3620
rect 13355 3595 13495 3600
rect 13355 3575 13405 3595
rect 13445 3575 13495 3595
rect 13535 3620 13675 3625
rect 13535 3600 13550 3620
rect 13570 3600 13640 3620
rect 13660 3600 13675 3620
rect 13535 3595 13675 3600
rect 13535 3575 13585 3595
rect 13625 3575 13675 3595
rect 13715 3620 13855 3625
rect 13715 3600 13730 3620
rect 13750 3600 13820 3620
rect 13840 3600 13855 3620
rect 13715 3595 13855 3600
rect 13715 3575 13765 3595
rect 13805 3575 13855 3595
rect 13895 3620 14035 3625
rect 13895 3600 13910 3620
rect 13930 3600 14000 3620
rect 14020 3600 14035 3620
rect 13895 3595 14035 3600
rect 13895 3575 13945 3595
rect 13985 3575 14035 3595
rect 14075 3620 14215 3625
rect 14075 3600 14090 3620
rect 14110 3600 14180 3620
rect 14200 3600 14215 3620
rect 14075 3595 14215 3600
rect 14075 3575 14125 3595
rect 14165 3575 14215 3595
rect 14255 3620 14395 3625
rect 14255 3600 14270 3620
rect 14290 3600 14360 3620
rect 14380 3600 14395 3620
rect 14255 3595 14395 3600
rect 14255 3575 14305 3595
rect 14345 3575 14395 3595
rect 14435 3620 14575 3625
rect 14435 3600 14450 3620
rect 14470 3600 14540 3620
rect 14560 3600 14575 3620
rect 14435 3595 14575 3600
rect 14435 3575 14485 3595
rect 14525 3575 14575 3595
rect 14615 3620 14755 3625
rect 14615 3600 14630 3620
rect 14650 3600 14720 3620
rect 14740 3600 14755 3620
rect 14615 3595 14755 3600
rect 14615 3575 14665 3595
rect 14705 3575 14755 3595
rect 14795 3620 14935 3625
rect 14795 3600 14810 3620
rect 14830 3600 14900 3620
rect 14920 3600 14935 3620
rect 14795 3595 14935 3600
rect 14795 3575 14845 3595
rect 14885 3575 14935 3595
rect 14975 3620 15115 3625
rect 14975 3600 14990 3620
rect 15010 3600 15080 3620
rect 15100 3600 15115 3620
rect 14975 3595 15115 3600
rect 14975 3575 15025 3595
rect 15065 3575 15115 3595
rect 15155 3620 15295 3625
rect 15155 3600 15170 3620
rect 15190 3600 15260 3620
rect 15280 3600 15295 3620
rect 15155 3595 15295 3600
rect 15155 3575 15205 3595
rect 15245 3575 15295 3595
rect 15335 3620 15475 3625
rect 15335 3600 15350 3620
rect 15370 3600 15440 3620
rect 15460 3600 15475 3620
rect 15335 3595 15475 3600
rect 15335 3575 15385 3595
rect 15425 3575 15475 3595
rect 15515 3620 15655 3625
rect 15515 3600 15530 3620
rect 15550 3600 15620 3620
rect 15640 3600 15655 3620
rect 15515 3595 15655 3600
rect 15515 3575 15565 3595
rect 15605 3575 15655 3595
rect 15695 3620 15835 3625
rect 15695 3600 15710 3620
rect 15730 3600 15800 3620
rect 15820 3600 15835 3620
rect 15695 3595 15835 3600
rect 15695 3575 15745 3595
rect 15785 3575 15835 3595
rect 15875 3620 16015 3625
rect 15875 3600 15890 3620
rect 15910 3600 15980 3620
rect 16000 3600 16015 3620
rect 15875 3595 16015 3600
rect 15875 3575 15925 3595
rect 15965 3575 16015 3595
rect 16055 3620 16195 3625
rect 16055 3600 16070 3620
rect 16090 3600 16160 3620
rect 16180 3600 16195 3620
rect 16055 3595 16195 3600
rect 16055 3575 16105 3595
rect 16145 3575 16195 3595
rect 16235 3620 16375 3625
rect 16235 3600 16250 3620
rect 16270 3600 16340 3620
rect 16360 3600 16375 3620
rect 16235 3595 16375 3600
rect 16235 3575 16285 3595
rect 16325 3575 16375 3595
rect 16415 3620 16555 3625
rect 16415 3600 16430 3620
rect 16450 3600 16520 3620
rect 16540 3600 16555 3620
rect 16415 3595 16555 3600
rect 16415 3575 16465 3595
rect 16505 3575 16555 3595
rect 16595 3620 16735 3625
rect 16595 3600 16610 3620
rect 16630 3600 16700 3620
rect 16720 3600 16735 3620
rect 16595 3595 16735 3600
rect 16595 3575 16645 3595
rect 16685 3575 16735 3595
rect 16775 3620 16915 3625
rect 16775 3600 16790 3620
rect 16810 3600 16880 3620
rect 16900 3600 16915 3620
rect 16775 3595 16915 3600
rect 16775 3575 16825 3595
rect 16865 3575 16915 3595
rect 16955 3620 17095 3625
rect 16955 3600 16970 3620
rect 16990 3600 17060 3620
rect 17080 3600 17095 3620
rect 16955 3595 17095 3600
rect 16955 3575 17005 3595
rect 17045 3575 17095 3595
rect 17135 3620 17275 3625
rect 17135 3600 17150 3620
rect 17170 3600 17240 3620
rect 17260 3600 17275 3620
rect 17135 3595 17275 3600
rect 17135 3575 17185 3595
rect 17225 3575 17275 3595
rect 17315 3620 17455 3625
rect 17315 3600 17330 3620
rect 17350 3600 17420 3620
rect 17440 3600 17455 3620
rect 17315 3595 17455 3600
rect 17315 3575 17365 3595
rect 17405 3575 17455 3595
rect 17495 3620 17635 3625
rect 17495 3600 17510 3620
rect 17530 3600 17600 3620
rect 17620 3600 17635 3620
rect 17495 3595 17635 3600
rect 17495 3575 17545 3595
rect 17585 3575 17635 3595
rect 17675 3620 17815 3625
rect 17675 3600 17690 3620
rect 17710 3600 17780 3620
rect 17800 3600 17815 3620
rect 17675 3595 17815 3600
rect 17675 3575 17725 3595
rect 17765 3575 17815 3595
rect 17855 3620 17995 3625
rect 17855 3600 17870 3620
rect 17890 3600 17960 3620
rect 17980 3600 17995 3620
rect 17855 3595 17995 3600
rect 17855 3575 17905 3595
rect 17945 3575 17995 3595
rect 18035 3620 18175 3625
rect 18035 3600 18050 3620
rect 18070 3600 18140 3620
rect 18160 3600 18175 3620
rect 18035 3595 18175 3600
rect 18035 3575 18085 3595
rect 18125 3575 18175 3595
rect 18215 3620 18355 3625
rect 18215 3600 18230 3620
rect 18250 3600 18320 3620
rect 18340 3600 18355 3620
rect 18215 3595 18355 3600
rect 18215 3575 18265 3595
rect 18305 3575 18355 3595
rect 18395 3620 18535 3625
rect 18395 3600 18410 3620
rect 18430 3600 18500 3620
rect 18520 3600 18535 3620
rect 18395 3595 18535 3600
rect 18395 3575 18445 3595
rect 18485 3575 18535 3595
rect 18575 3620 18715 3625
rect 18575 3600 18590 3620
rect 18610 3600 18680 3620
rect 18700 3600 18715 3620
rect 18575 3595 18715 3600
rect 18575 3575 18625 3595
rect 18665 3575 18715 3595
rect 18755 3620 18895 3625
rect 18755 3600 18770 3620
rect 18790 3600 18860 3620
rect 18880 3600 18895 3620
rect 18755 3595 18895 3600
rect 18755 3575 18805 3595
rect 18845 3575 18895 3595
rect 18935 3620 19075 3625
rect 18935 3600 18950 3620
rect 18970 3600 19040 3620
rect 19060 3600 19075 3620
rect 18935 3595 19075 3600
rect 18935 3575 18985 3595
rect 19025 3575 19075 3595
rect 19115 3620 19255 3625
rect 19115 3600 19130 3620
rect 19150 3600 19220 3620
rect 19240 3600 19255 3620
rect 19115 3595 19255 3600
rect 19115 3575 19165 3595
rect 19205 3575 19255 3595
rect 19295 3620 19435 3625
rect 19295 3600 19310 3620
rect 19330 3600 19400 3620
rect 19420 3600 19435 3620
rect 19295 3595 19435 3600
rect 19295 3575 19345 3595
rect 19385 3575 19435 3595
rect 19475 3620 19615 3625
rect 19475 3600 19490 3620
rect 19510 3600 19580 3620
rect 19600 3600 19615 3620
rect 19475 3595 19615 3600
rect 19475 3575 19525 3595
rect 19565 3575 19615 3595
rect 19655 3620 19795 3625
rect 19655 3600 19670 3620
rect 19690 3600 19760 3620
rect 19780 3600 19795 3620
rect 19655 3595 19795 3600
rect 19655 3575 19705 3595
rect 19745 3575 19795 3595
rect 19835 3620 19975 3625
rect 19835 3600 19850 3620
rect 19870 3600 19940 3620
rect 19960 3600 19975 3620
rect 19835 3595 19975 3600
rect 19835 3575 19885 3595
rect 19925 3575 19975 3595
rect 20015 3620 20155 3625
rect 20015 3600 20030 3620
rect 20050 3600 20120 3620
rect 20140 3600 20155 3620
rect 20015 3595 20155 3600
rect 20015 3575 20065 3595
rect 20105 3575 20155 3595
rect 20195 3620 20335 3625
rect 20195 3600 20210 3620
rect 20230 3600 20300 3620
rect 20320 3600 20335 3620
rect 20195 3595 20335 3600
rect 20195 3575 20245 3595
rect 20285 3575 20335 3595
rect 20375 3620 20515 3625
rect 20375 3600 20390 3620
rect 20410 3600 20480 3620
rect 20500 3600 20515 3620
rect 20375 3595 20515 3600
rect 20375 3575 20425 3595
rect 20465 3575 20515 3595
rect 20555 3620 20695 3625
rect 20555 3600 20570 3620
rect 20590 3600 20660 3620
rect 20680 3600 20695 3620
rect 20555 3595 20695 3600
rect 20555 3575 20605 3595
rect 20645 3575 20695 3595
rect 9215 3460 9265 3475
rect 9305 3460 9355 3475
rect 9395 3460 9445 3475
rect 9485 3460 9535 3475
rect 9575 3460 9625 3475
rect 9665 3460 9715 3475
rect 9755 3460 9805 3475
rect 9845 3460 9895 3475
rect 9935 3460 9985 3475
rect 10025 3460 10075 3475
rect 10115 3460 10165 3475
rect 10205 3460 10255 3475
rect 10295 3460 10345 3475
rect 10385 3460 10435 3475
rect 10475 3460 10525 3475
rect 10565 3460 10615 3475
rect 10655 3460 10705 3475
rect 10745 3460 10795 3475
rect 10835 3460 10885 3475
rect 10925 3460 10975 3475
rect 11015 3460 11065 3475
rect 11105 3460 11155 3475
rect 11195 3460 11245 3475
rect 11285 3460 11335 3475
rect 11375 3460 11425 3475
rect 11465 3460 11515 3475
rect 11555 3460 11605 3475
rect 11645 3460 11695 3475
rect 11735 3460 11785 3475
rect 11825 3460 11875 3475
rect 11915 3460 11965 3475
rect 12005 3460 12055 3475
rect 12095 3460 12145 3475
rect 12185 3460 12235 3475
rect 12275 3460 12325 3475
rect 12365 3460 12415 3475
rect 12455 3460 12505 3475
rect 12545 3460 12595 3475
rect 12635 3460 12685 3475
rect 12725 3460 12775 3475
rect 12815 3460 12865 3475
rect 12905 3460 12955 3475
rect 12995 3460 13045 3475
rect 13085 3460 13135 3475
rect 13175 3460 13225 3475
rect 13265 3460 13315 3475
rect 13355 3460 13405 3475
rect 13445 3460 13495 3475
rect 13535 3460 13585 3475
rect 13625 3460 13675 3475
rect 13715 3460 13765 3475
rect 13805 3460 13855 3475
rect 13895 3460 13945 3475
rect 13985 3460 14035 3475
rect 14075 3460 14125 3475
rect 14165 3460 14215 3475
rect 14255 3460 14305 3475
rect 14345 3460 14395 3475
rect 14435 3460 14485 3475
rect 14525 3460 14575 3475
rect 14615 3460 14665 3475
rect 14705 3460 14755 3475
rect 14795 3460 14845 3475
rect 14885 3460 14935 3475
rect 14975 3460 15025 3475
rect 15065 3460 15115 3475
rect 15155 3460 15205 3475
rect 15245 3460 15295 3475
rect 15335 3460 15385 3475
rect 15425 3460 15475 3475
rect 15515 3460 15565 3475
rect 15605 3460 15655 3475
rect 15695 3460 15745 3475
rect 15785 3460 15835 3475
rect 15875 3460 15925 3475
rect 15965 3460 16015 3475
rect 16055 3460 16105 3475
rect 16145 3460 16195 3475
rect 16235 3460 16285 3475
rect 16325 3460 16375 3475
rect 16415 3460 16465 3475
rect 16505 3460 16555 3475
rect 16595 3460 16645 3475
rect 16685 3460 16735 3475
rect 16775 3460 16825 3475
rect 16865 3460 16915 3475
rect 16955 3460 17005 3475
rect 17045 3460 17095 3475
rect 17135 3460 17185 3475
rect 17225 3460 17275 3475
rect 17315 3460 17365 3475
rect 17405 3460 17455 3475
rect 17495 3460 17545 3475
rect 17585 3460 17635 3475
rect 17675 3460 17725 3475
rect 17765 3460 17815 3475
rect 17855 3460 17905 3475
rect 17945 3460 17995 3475
rect 18035 3460 18085 3475
rect 18125 3460 18175 3475
rect 18215 3460 18265 3475
rect 18305 3460 18355 3475
rect 18395 3460 18445 3475
rect 18485 3460 18535 3475
rect 18575 3460 18625 3475
rect 18665 3460 18715 3475
rect 18755 3460 18805 3475
rect 18845 3460 18895 3475
rect 18935 3460 18985 3475
rect 19025 3460 19075 3475
rect 19115 3460 19165 3475
rect 19205 3460 19255 3475
rect 19295 3460 19345 3475
rect 19385 3460 19435 3475
rect 19475 3460 19525 3475
rect 19565 3460 19615 3475
rect 19655 3460 19705 3475
rect 19745 3460 19795 3475
rect 19835 3460 19885 3475
rect 19925 3460 19975 3475
rect 20015 3460 20065 3475
rect 20105 3460 20155 3475
rect 20195 3460 20245 3475
rect 20285 3460 20335 3475
rect 20375 3460 20425 3475
rect 20465 3460 20515 3475
rect 20555 3460 20605 3475
rect 20645 3460 20695 3475
<< polycont >>
rect 9230 4170 9250 4190
rect 9320 4170 9340 4190
rect 9410 4170 9430 4190
rect 9500 4170 9520 4190
rect 9590 4170 9610 4190
rect 9680 4170 9700 4190
rect 9770 4170 9790 4190
rect 9860 4170 9880 4190
rect 9950 4170 9970 4190
rect 10040 4170 10060 4190
rect 10130 4170 10150 4190
rect 10220 4170 10240 4190
rect 10310 4170 10330 4190
rect 10400 4170 10420 4190
rect 10490 4170 10510 4190
rect 10580 4170 10600 4190
rect 10670 4170 10690 4190
rect 10760 4170 10780 4190
rect 10850 4170 10870 4190
rect 10940 4170 10960 4190
rect 11030 4170 11050 4190
rect 11120 4170 11140 4190
rect 11210 4170 11230 4190
rect 11300 4170 11320 4190
rect 11390 4170 11410 4190
rect 11480 4170 11500 4190
rect 11570 4170 11590 4190
rect 11660 4170 11680 4190
rect 11750 4170 11770 4190
rect 11840 4170 11860 4190
rect 11930 4170 11950 4190
rect 12020 4170 12040 4190
rect 12110 4170 12130 4190
rect 12200 4170 12220 4190
rect 12290 4170 12310 4190
rect 12380 4170 12400 4190
rect 12470 4170 12490 4190
rect 12560 4170 12580 4190
rect 12650 4170 12670 4190
rect 12740 4170 12760 4190
rect 12830 4170 12850 4190
rect 12920 4170 12940 4190
rect 13010 4170 13030 4190
rect 13100 4170 13120 4190
rect 13190 4170 13210 4190
rect 13280 4170 13300 4190
rect 13370 4170 13390 4190
rect 13460 4170 13480 4190
rect 13550 4170 13570 4190
rect 13640 4170 13660 4190
rect 13730 4170 13750 4190
rect 13820 4170 13840 4190
rect 13910 4170 13930 4190
rect 14000 4170 14020 4190
rect 14090 4170 14110 4190
rect 14180 4170 14200 4190
rect 14270 4170 14290 4190
rect 14360 4170 14380 4190
rect 14450 4170 14470 4190
rect 14540 4170 14560 4190
rect 14630 4170 14650 4190
rect 14720 4170 14740 4190
rect 14810 4170 14830 4190
rect 14900 4170 14920 4190
rect 14990 4170 15010 4190
rect 15080 4170 15100 4190
rect 15170 4170 15190 4190
rect 15260 4170 15280 4190
rect 15350 4170 15370 4190
rect 15440 4170 15460 4190
rect 15530 4170 15550 4190
rect 15620 4170 15640 4190
rect 15710 4170 15730 4190
rect 15800 4170 15820 4190
rect 15890 4170 15910 4190
rect 15980 4170 16000 4190
rect 16070 4170 16090 4190
rect 16160 4170 16180 4190
rect 16250 4170 16270 4190
rect 16340 4170 16360 4190
rect 16430 4170 16450 4190
rect 16520 4170 16540 4190
rect 16610 4170 16630 4190
rect 16700 4170 16720 4190
rect 16790 4170 16810 4190
rect 16880 4170 16900 4190
rect 16970 4170 16990 4190
rect 17060 4170 17080 4190
rect 17150 4170 17170 4190
rect 17240 4170 17260 4190
rect 17330 4170 17350 4190
rect 17420 4170 17440 4190
rect 17510 4170 17530 4190
rect 17600 4170 17620 4190
rect 17690 4170 17710 4190
rect 17780 4170 17800 4190
rect 17870 4170 17890 4190
rect 17960 4170 17980 4190
rect 18050 4170 18070 4190
rect 18140 4170 18160 4190
rect 18230 4170 18250 4190
rect 18320 4170 18340 4190
rect 18410 4170 18430 4190
rect 18500 4170 18520 4190
rect 18590 4170 18610 4190
rect 18680 4170 18700 4190
rect 18770 4170 18790 4190
rect 18860 4170 18880 4190
rect 18950 4170 18970 4190
rect 19040 4170 19060 4190
rect 19130 4170 19150 4190
rect 19220 4170 19240 4190
rect 19310 4170 19330 4190
rect 19400 4170 19420 4190
rect 19490 4170 19510 4190
rect 19580 4170 19600 4190
rect 19670 4170 19690 4190
rect 19760 4170 19780 4190
rect 19850 4170 19870 4190
rect 19940 4170 19960 4190
rect 20030 4170 20050 4190
rect 20120 4170 20140 4190
rect 20210 4170 20230 4190
rect 20300 4170 20320 4190
rect 20390 4170 20410 4190
rect 20480 4170 20500 4190
rect 20570 4170 20590 4190
rect 20660 4170 20680 4190
rect 9230 3600 9250 3620
rect 9320 3600 9340 3620
rect 9410 3600 9430 3620
rect 9500 3600 9520 3620
rect 9590 3600 9610 3620
rect 9680 3600 9700 3620
rect 9770 3600 9790 3620
rect 9860 3600 9880 3620
rect 9950 3600 9970 3620
rect 10040 3600 10060 3620
rect 10130 3600 10150 3620
rect 10220 3600 10240 3620
rect 10310 3600 10330 3620
rect 10400 3600 10420 3620
rect 10490 3600 10510 3620
rect 10580 3600 10600 3620
rect 10670 3600 10690 3620
rect 10760 3600 10780 3620
rect 10850 3600 10870 3620
rect 10940 3600 10960 3620
rect 11030 3600 11050 3620
rect 11120 3600 11140 3620
rect 11210 3600 11230 3620
rect 11300 3600 11320 3620
rect 11390 3600 11410 3620
rect 11480 3600 11500 3620
rect 11570 3600 11590 3620
rect 11660 3600 11680 3620
rect 11750 3600 11770 3620
rect 11840 3600 11860 3620
rect 11930 3600 11950 3620
rect 12020 3600 12040 3620
rect 12110 3600 12130 3620
rect 12200 3600 12220 3620
rect 12290 3600 12310 3620
rect 12380 3600 12400 3620
rect 12470 3600 12490 3620
rect 12560 3600 12580 3620
rect 12650 3600 12670 3620
rect 12740 3600 12760 3620
rect 12830 3600 12850 3620
rect 12920 3600 12940 3620
rect 13010 3600 13030 3620
rect 13100 3600 13120 3620
rect 13190 3600 13210 3620
rect 13280 3600 13300 3620
rect 13370 3600 13390 3620
rect 13460 3600 13480 3620
rect 13550 3600 13570 3620
rect 13640 3600 13660 3620
rect 13730 3600 13750 3620
rect 13820 3600 13840 3620
rect 13910 3600 13930 3620
rect 14000 3600 14020 3620
rect 14090 3600 14110 3620
rect 14180 3600 14200 3620
rect 14270 3600 14290 3620
rect 14360 3600 14380 3620
rect 14450 3600 14470 3620
rect 14540 3600 14560 3620
rect 14630 3600 14650 3620
rect 14720 3600 14740 3620
rect 14810 3600 14830 3620
rect 14900 3600 14920 3620
rect 14990 3600 15010 3620
rect 15080 3600 15100 3620
rect 15170 3600 15190 3620
rect 15260 3600 15280 3620
rect 15350 3600 15370 3620
rect 15440 3600 15460 3620
rect 15530 3600 15550 3620
rect 15620 3600 15640 3620
rect 15710 3600 15730 3620
rect 15800 3600 15820 3620
rect 15890 3600 15910 3620
rect 15980 3600 16000 3620
rect 16070 3600 16090 3620
rect 16160 3600 16180 3620
rect 16250 3600 16270 3620
rect 16340 3600 16360 3620
rect 16430 3600 16450 3620
rect 16520 3600 16540 3620
rect 16610 3600 16630 3620
rect 16700 3600 16720 3620
rect 16790 3600 16810 3620
rect 16880 3600 16900 3620
rect 16970 3600 16990 3620
rect 17060 3600 17080 3620
rect 17150 3600 17170 3620
rect 17240 3600 17260 3620
rect 17330 3600 17350 3620
rect 17420 3600 17440 3620
rect 17510 3600 17530 3620
rect 17600 3600 17620 3620
rect 17690 3600 17710 3620
rect 17780 3600 17800 3620
rect 17870 3600 17890 3620
rect 17960 3600 17980 3620
rect 18050 3600 18070 3620
rect 18140 3600 18160 3620
rect 18230 3600 18250 3620
rect 18320 3600 18340 3620
rect 18410 3600 18430 3620
rect 18500 3600 18520 3620
rect 18590 3600 18610 3620
rect 18680 3600 18700 3620
rect 18770 3600 18790 3620
rect 18860 3600 18880 3620
rect 18950 3600 18970 3620
rect 19040 3600 19060 3620
rect 19130 3600 19150 3620
rect 19220 3600 19240 3620
rect 19310 3600 19330 3620
rect 19400 3600 19420 3620
rect 19490 3600 19510 3620
rect 19580 3600 19600 3620
rect 19670 3600 19690 3620
rect 19760 3600 19780 3620
rect 19850 3600 19870 3620
rect 19940 3600 19960 3620
rect 20030 3600 20050 3620
rect 20120 3600 20140 3620
rect 20210 3600 20230 3620
rect 20300 3600 20320 3620
rect 20390 3600 20410 3620
rect 20480 3600 20500 3620
rect 20570 3600 20590 3620
rect 20660 3600 20680 3620
<< locali >>
rect 9050 4065 9070 4375
rect 9125 4345 9185 4365
rect 9205 4345 9230 4365
rect 9250 4345 9320 4365
rect 9340 4345 9410 4365
rect 9430 4345 9500 4365
rect 9520 4345 9590 4365
rect 9610 4345 9680 4365
rect 9700 4345 9770 4365
rect 9790 4345 9860 4365
rect 9880 4345 9905 4365
rect 9925 4345 9950 4365
rect 9970 4345 10040 4365
rect 10060 4345 10085 4365
rect 10105 4345 10130 4365
rect 10150 4345 10220 4365
rect 10240 4345 10265 4365
rect 10285 4345 10310 4365
rect 10330 4345 10400 4365
rect 10420 4345 10445 4365
rect 10465 4345 10490 4365
rect 10510 4345 10580 4365
rect 10600 4345 10625 4365
rect 10645 4345 10670 4365
rect 10690 4345 10760 4365
rect 10780 4345 10805 4365
rect 10825 4345 10850 4365
rect 10870 4345 10940 4365
rect 10960 4345 10985 4365
rect 11005 4345 11030 4365
rect 11050 4345 11120 4365
rect 11140 4345 11165 4365
rect 11185 4345 11210 4365
rect 11230 4345 11300 4365
rect 11320 4345 11345 4365
rect 11365 4345 11390 4365
rect 11410 4345 11480 4365
rect 11500 4345 11525 4365
rect 11545 4345 11570 4365
rect 11590 4345 11660 4365
rect 11680 4345 11705 4365
rect 11725 4345 11750 4365
rect 11770 4345 11840 4365
rect 11860 4345 11885 4365
rect 11905 4345 11930 4365
rect 11950 4345 12020 4365
rect 12040 4345 12065 4365
rect 12085 4345 12110 4365
rect 12130 4345 12200 4365
rect 12220 4345 12245 4365
rect 12265 4345 12290 4365
rect 12310 4345 12380 4365
rect 12400 4345 12425 4365
rect 12445 4345 12470 4365
rect 12490 4345 12560 4365
rect 12580 4345 12605 4365
rect 12625 4345 12650 4365
rect 12670 4345 12740 4365
rect 12760 4345 12785 4365
rect 12805 4345 12830 4365
rect 12850 4345 12920 4365
rect 12940 4345 12965 4365
rect 12985 4345 13010 4365
rect 13030 4345 13100 4365
rect 13120 4345 13145 4365
rect 13165 4345 13190 4365
rect 13210 4345 13280 4365
rect 13300 4345 13325 4365
rect 13345 4345 13370 4365
rect 13390 4345 13460 4365
rect 13480 4345 13505 4365
rect 13525 4345 13550 4365
rect 13570 4345 13640 4365
rect 13660 4345 13685 4365
rect 13705 4345 13730 4365
rect 13750 4345 13820 4365
rect 13840 4345 13865 4365
rect 13885 4345 13910 4365
rect 13930 4345 14000 4365
rect 14020 4345 14045 4365
rect 14065 4345 14090 4365
rect 14110 4345 14180 4365
rect 14200 4345 14225 4365
rect 14245 4345 14270 4365
rect 14290 4345 14360 4365
rect 14380 4345 14405 4365
rect 14425 4345 14450 4365
rect 14470 4345 14540 4365
rect 14560 4345 14585 4365
rect 14605 4345 14630 4365
rect 14650 4345 14720 4365
rect 14740 4345 14765 4365
rect 14785 4345 14810 4365
rect 14830 4345 14900 4365
rect 14920 4345 14945 4365
rect 14965 4345 14990 4365
rect 15010 4345 15080 4365
rect 15100 4345 15125 4365
rect 15145 4345 15170 4365
rect 15190 4345 15260 4365
rect 15280 4345 15305 4365
rect 15325 4345 15350 4365
rect 15370 4345 15440 4365
rect 15460 4345 15485 4365
rect 15505 4345 15530 4365
rect 15550 4345 15620 4365
rect 15640 4345 15665 4365
rect 15685 4345 15710 4365
rect 15730 4345 15800 4365
rect 15820 4345 15845 4365
rect 15865 4345 15890 4365
rect 15910 4345 15980 4365
rect 16000 4345 16025 4365
rect 16045 4345 16070 4365
rect 16090 4345 16160 4365
rect 16180 4345 16205 4365
rect 16225 4345 16250 4365
rect 16270 4345 16340 4365
rect 16360 4345 16385 4365
rect 16405 4345 16430 4365
rect 16450 4345 16520 4365
rect 16540 4345 16565 4365
rect 16585 4345 16610 4365
rect 16630 4345 16700 4365
rect 16720 4345 16745 4365
rect 16765 4345 16790 4365
rect 16810 4345 16880 4365
rect 16900 4345 16925 4365
rect 16945 4345 16970 4365
rect 16990 4345 17060 4365
rect 17080 4345 17105 4365
rect 17125 4345 17150 4365
rect 17170 4345 17240 4365
rect 17260 4345 17285 4365
rect 17305 4345 17330 4365
rect 17350 4345 17420 4365
rect 17440 4345 17465 4365
rect 17485 4345 17510 4365
rect 17530 4345 17600 4365
rect 17620 4345 17645 4365
rect 17665 4345 17690 4365
rect 17710 4345 17780 4365
rect 17800 4345 17825 4365
rect 17845 4345 17870 4365
rect 17890 4345 17960 4365
rect 17980 4345 18005 4365
rect 18025 4345 18050 4365
rect 18070 4345 18140 4365
rect 18160 4345 18185 4365
rect 18205 4345 18230 4365
rect 18250 4345 18320 4365
rect 18340 4345 18365 4365
rect 18385 4345 18410 4365
rect 18430 4345 18500 4365
rect 18520 4345 18545 4365
rect 18565 4345 18590 4365
rect 18610 4345 18680 4365
rect 18700 4345 18725 4365
rect 18745 4345 18770 4365
rect 18790 4345 18860 4365
rect 18880 4345 18905 4365
rect 18925 4345 18950 4365
rect 18970 4345 19040 4365
rect 19060 4345 19085 4365
rect 19105 4345 19130 4365
rect 19150 4345 19220 4365
rect 19240 4345 19265 4365
rect 19285 4345 19310 4365
rect 19330 4345 19400 4365
rect 19420 4345 19445 4365
rect 19465 4345 19490 4365
rect 19510 4345 19580 4365
rect 19600 4345 19625 4365
rect 19645 4345 19670 4365
rect 19690 4345 19760 4365
rect 19780 4345 19805 4365
rect 19825 4345 19850 4365
rect 19870 4345 19940 4365
rect 19960 4345 19985 4365
rect 20005 4345 20030 4365
rect 20050 4345 20120 4365
rect 20140 4345 20210 4365
rect 20230 4345 20300 4365
rect 20320 4345 20390 4365
rect 20410 4345 20480 4365
rect 20500 4345 20570 4365
rect 20590 4345 20660 4365
rect 20680 4345 20705 4365
rect 20725 4345 20785 4365
rect 9125 4145 9145 4345
rect 9185 4305 9205 4315
rect 9185 4215 9205 4225
rect 9275 4305 9295 4315
rect 9275 4215 9295 4225
rect 9365 4305 9385 4315
rect 9365 4215 9385 4225
rect 9455 4305 9475 4315
rect 9455 4190 9475 4225
rect 9545 4305 9565 4315
rect 9545 4215 9565 4225
rect 9635 4305 9655 4315
rect 9635 4190 9655 4225
rect 9725 4305 9745 4315
rect 9725 4215 9745 4225
rect 9815 4305 9835 4315
rect 9815 4215 9835 4225
rect 9905 4305 9925 4315
rect 9905 4215 9925 4225
rect 9995 4305 10015 4315
rect 9995 4215 10015 4225
rect 10085 4305 10105 4315
rect 10085 4215 10105 4225
rect 10175 4305 10195 4315
rect 10175 4215 10195 4225
rect 10265 4305 10285 4315
rect 10265 4215 10285 4225
rect 10355 4305 10375 4315
rect 10355 4215 10375 4225
rect 10445 4305 10465 4315
rect 10445 4215 10465 4225
rect 10535 4305 10555 4315
rect 10535 4215 10555 4225
rect 10625 4305 10645 4315
rect 10625 4215 10645 4225
rect 10715 4305 10735 4315
rect 10715 4215 10735 4225
rect 10805 4305 10825 4315
rect 10805 4215 10825 4225
rect 10895 4305 10915 4315
rect 10895 4215 10915 4225
rect 10985 4305 11005 4315
rect 10985 4215 11005 4225
rect 11075 4305 11095 4315
rect 11075 4215 11095 4225
rect 11165 4305 11185 4315
rect 11165 4215 11185 4225
rect 11255 4305 11275 4315
rect 11255 4215 11275 4225
rect 11345 4305 11365 4315
rect 11345 4215 11365 4225
rect 11435 4305 11455 4315
rect 11435 4215 11455 4225
rect 11525 4305 11545 4315
rect 11525 4215 11545 4225
rect 11615 4305 11635 4315
rect 11615 4215 11635 4225
rect 11705 4305 11725 4315
rect 11705 4215 11725 4225
rect 11795 4305 11815 4315
rect 11795 4215 11815 4225
rect 11885 4305 11905 4315
rect 11885 4215 11905 4225
rect 11975 4305 11995 4315
rect 11975 4215 11995 4225
rect 12065 4305 12085 4315
rect 12065 4215 12085 4225
rect 12155 4305 12175 4315
rect 12155 4215 12175 4225
rect 12245 4305 12265 4315
rect 12245 4215 12265 4225
rect 12335 4305 12355 4315
rect 12335 4215 12355 4225
rect 12425 4305 12445 4315
rect 12425 4215 12445 4225
rect 12515 4305 12535 4315
rect 12515 4215 12535 4225
rect 12605 4305 12625 4315
rect 12605 4215 12625 4225
rect 12695 4305 12715 4315
rect 12695 4215 12715 4225
rect 12785 4305 12805 4315
rect 12785 4215 12805 4225
rect 12875 4305 12895 4315
rect 12875 4215 12895 4225
rect 12965 4305 12985 4315
rect 12965 4215 12985 4225
rect 13055 4305 13075 4315
rect 13055 4215 13075 4225
rect 13145 4305 13165 4315
rect 13145 4215 13165 4225
rect 13235 4305 13255 4315
rect 13235 4215 13255 4225
rect 13325 4305 13345 4315
rect 13325 4215 13345 4225
rect 13415 4305 13435 4315
rect 13415 4215 13435 4225
rect 13505 4305 13525 4315
rect 13505 4215 13525 4225
rect 13595 4305 13615 4315
rect 13595 4215 13615 4225
rect 13685 4305 13705 4315
rect 13685 4215 13705 4225
rect 13775 4305 13795 4315
rect 13775 4215 13795 4225
rect 13865 4305 13885 4315
rect 13865 4215 13885 4225
rect 13955 4305 13975 4315
rect 13955 4215 13975 4225
rect 14045 4305 14065 4315
rect 14045 4215 14065 4225
rect 14135 4305 14155 4315
rect 14135 4215 14155 4225
rect 14225 4305 14245 4315
rect 14225 4215 14245 4225
rect 14315 4305 14335 4315
rect 14315 4215 14335 4225
rect 14405 4305 14425 4315
rect 14405 4215 14425 4225
rect 14495 4305 14515 4315
rect 14495 4215 14515 4225
rect 14585 4305 14605 4315
rect 14585 4215 14605 4225
rect 14675 4305 14695 4315
rect 14675 4215 14695 4225
rect 14765 4305 14785 4315
rect 14765 4215 14785 4225
rect 14855 4305 14875 4315
rect 14855 4215 14875 4225
rect 14945 4305 14965 4315
rect 14945 4215 14965 4225
rect 15035 4305 15055 4315
rect 15035 4215 15055 4225
rect 15125 4305 15145 4315
rect 15125 4215 15145 4225
rect 15215 4305 15235 4315
rect 15215 4215 15235 4225
rect 15305 4305 15325 4315
rect 15305 4215 15325 4225
rect 15395 4305 15415 4315
rect 15395 4215 15415 4225
rect 15485 4305 15505 4315
rect 15485 4215 15505 4225
rect 15575 4305 15595 4315
rect 15575 4215 15595 4225
rect 15665 4305 15685 4315
rect 15665 4215 15685 4225
rect 15755 4305 15775 4315
rect 15755 4215 15775 4225
rect 15845 4305 15865 4315
rect 15845 4215 15865 4225
rect 15935 4305 15955 4315
rect 15935 4215 15955 4225
rect 16025 4305 16045 4315
rect 16025 4215 16045 4225
rect 16115 4305 16135 4315
rect 16115 4215 16135 4225
rect 16205 4305 16225 4315
rect 16205 4215 16225 4225
rect 16295 4305 16315 4315
rect 16295 4215 16315 4225
rect 16385 4305 16405 4315
rect 16385 4215 16405 4225
rect 16475 4305 16495 4315
rect 16475 4215 16495 4225
rect 16565 4305 16585 4315
rect 16565 4215 16585 4225
rect 16655 4305 16675 4315
rect 16655 4215 16675 4225
rect 16745 4305 16765 4315
rect 16745 4215 16765 4225
rect 16835 4305 16855 4315
rect 16835 4215 16855 4225
rect 16925 4305 16945 4315
rect 16925 4215 16945 4225
rect 17015 4305 17035 4315
rect 17015 4215 17035 4225
rect 17105 4305 17125 4315
rect 17105 4215 17125 4225
rect 17195 4305 17215 4315
rect 17195 4215 17215 4225
rect 17285 4305 17305 4315
rect 17285 4215 17305 4225
rect 17375 4305 17395 4315
rect 17375 4215 17395 4225
rect 17465 4305 17485 4315
rect 17465 4215 17485 4225
rect 17555 4305 17575 4315
rect 17555 4215 17575 4225
rect 17645 4305 17665 4315
rect 17645 4215 17665 4225
rect 17735 4305 17755 4315
rect 17735 4215 17755 4225
rect 17825 4305 17845 4315
rect 17825 4215 17845 4225
rect 17915 4305 17935 4315
rect 17915 4215 17935 4225
rect 18005 4305 18025 4315
rect 18005 4215 18025 4225
rect 18095 4305 18115 4315
rect 18095 4215 18115 4225
rect 18185 4305 18205 4315
rect 18185 4215 18205 4225
rect 18275 4305 18295 4315
rect 18275 4215 18295 4225
rect 18365 4305 18385 4315
rect 18365 4215 18385 4225
rect 18455 4305 18475 4315
rect 18455 4215 18475 4225
rect 18545 4305 18565 4315
rect 18545 4215 18565 4225
rect 18635 4305 18655 4315
rect 18635 4215 18655 4225
rect 18725 4305 18745 4315
rect 18725 4215 18745 4225
rect 18815 4305 18835 4315
rect 18815 4215 18835 4225
rect 18905 4305 18925 4315
rect 18905 4215 18925 4225
rect 18995 4305 19015 4315
rect 18995 4215 19015 4225
rect 19085 4305 19105 4315
rect 19085 4215 19105 4225
rect 19175 4305 19195 4315
rect 19175 4215 19195 4225
rect 19265 4305 19285 4315
rect 19265 4215 19285 4225
rect 19355 4305 19375 4315
rect 19355 4215 19375 4225
rect 19445 4305 19465 4315
rect 19445 4215 19465 4225
rect 19535 4305 19555 4315
rect 19535 4215 19555 4225
rect 19625 4305 19645 4315
rect 19625 4215 19645 4225
rect 19715 4305 19735 4315
rect 19715 4215 19735 4225
rect 19805 4305 19825 4315
rect 19805 4215 19825 4225
rect 19895 4305 19915 4315
rect 19895 4215 19915 4225
rect 19985 4305 20005 4315
rect 19985 4215 20005 4225
rect 20075 4305 20095 4315
rect 20075 4215 20095 4225
rect 20165 4305 20185 4315
rect 20165 4215 20185 4225
rect 20255 4305 20275 4315
rect 20255 4190 20275 4225
rect 20345 4305 20365 4315
rect 20345 4215 20365 4225
rect 20435 4305 20455 4315
rect 20435 4190 20455 4225
rect 20525 4305 20545 4315
rect 20525 4215 20545 4225
rect 20615 4305 20635 4315
rect 20615 4215 20635 4225
rect 20705 4305 20725 4315
rect 20705 4215 20725 4225
rect 9220 4170 9230 4190
rect 9250 4170 9320 4190
rect 9340 4170 9410 4190
rect 9430 4170 9500 4190
rect 9520 4170 9590 4190
rect 9610 4170 9680 4190
rect 9700 4170 9770 4190
rect 9790 4170 9860 4190
rect 9880 4170 9895 4190
rect 9940 4170 9950 4190
rect 9970 4170 10040 4190
rect 10060 4170 10070 4190
rect 10120 4170 10130 4190
rect 10150 4170 10220 4190
rect 10240 4170 10250 4190
rect 10300 4170 10310 4190
rect 10330 4170 10400 4190
rect 10420 4170 10430 4190
rect 10480 4170 10490 4190
rect 10510 4170 10580 4190
rect 10600 4170 10610 4190
rect 10660 4170 10670 4190
rect 10690 4170 10760 4190
rect 10780 4170 10790 4190
rect 10840 4170 10850 4190
rect 10870 4170 10940 4190
rect 10960 4170 10970 4190
rect 11020 4170 11030 4190
rect 11050 4170 11120 4190
rect 11140 4170 11150 4190
rect 11200 4170 11210 4190
rect 11230 4170 11300 4190
rect 11320 4170 11330 4190
rect 11380 4170 11390 4190
rect 11410 4170 11480 4190
rect 11500 4170 11510 4190
rect 11560 4170 11570 4190
rect 11590 4170 11660 4190
rect 11680 4170 11690 4190
rect 11740 4170 11750 4190
rect 11770 4170 11840 4190
rect 11860 4170 11870 4190
rect 11920 4170 11930 4190
rect 11950 4170 12020 4190
rect 12040 4170 12050 4190
rect 12100 4170 12110 4190
rect 12130 4170 12200 4190
rect 12220 4170 12230 4190
rect 12280 4170 12290 4190
rect 12310 4170 12380 4190
rect 12400 4170 12410 4190
rect 12460 4170 12470 4190
rect 12490 4170 12560 4190
rect 12580 4170 12590 4190
rect 12640 4170 12650 4190
rect 12670 4170 12740 4190
rect 12760 4170 12770 4190
rect 12820 4170 12830 4190
rect 12850 4170 12920 4190
rect 12940 4170 12950 4190
rect 13000 4170 13010 4190
rect 13030 4170 13100 4190
rect 13120 4170 13130 4190
rect 13180 4170 13190 4190
rect 13210 4170 13280 4190
rect 13300 4170 13310 4190
rect 13360 4170 13370 4190
rect 13390 4170 13460 4190
rect 13480 4170 13490 4190
rect 13540 4170 13550 4190
rect 13570 4170 13640 4190
rect 13660 4170 13670 4190
rect 13720 4170 13730 4190
rect 13750 4170 13820 4190
rect 13840 4170 13850 4190
rect 13900 4170 13910 4190
rect 13930 4170 14000 4190
rect 14020 4170 14030 4190
rect 14080 4170 14090 4190
rect 14110 4170 14180 4190
rect 14200 4170 14210 4190
rect 14260 4170 14270 4190
rect 14290 4170 14360 4190
rect 14380 4170 14390 4190
rect 14440 4170 14450 4190
rect 14470 4170 14540 4190
rect 14560 4170 14570 4190
rect 14620 4170 14630 4190
rect 14650 4170 14720 4190
rect 14740 4170 14750 4190
rect 14800 4170 14810 4190
rect 14830 4170 14900 4190
rect 14920 4170 14930 4190
rect 14980 4170 14990 4190
rect 15010 4170 15080 4190
rect 15100 4170 15110 4190
rect 15160 4170 15170 4190
rect 15190 4170 15260 4190
rect 15280 4170 15290 4190
rect 15340 4170 15350 4190
rect 15370 4170 15440 4190
rect 15460 4170 15470 4190
rect 15520 4170 15530 4190
rect 15550 4170 15620 4190
rect 15640 4170 15650 4190
rect 15700 4170 15710 4190
rect 15730 4170 15800 4190
rect 15820 4170 15830 4190
rect 15880 4170 15890 4190
rect 15910 4170 15980 4190
rect 16000 4170 16010 4190
rect 16060 4170 16070 4190
rect 16090 4170 16160 4190
rect 16180 4170 16190 4190
rect 16240 4170 16250 4190
rect 16270 4170 16340 4190
rect 16360 4170 16370 4190
rect 16420 4170 16430 4190
rect 16450 4170 16520 4190
rect 16540 4170 16550 4190
rect 16600 4170 16610 4190
rect 16630 4170 16700 4190
rect 16720 4170 16730 4190
rect 16780 4170 16790 4190
rect 16810 4170 16880 4190
rect 16900 4170 16910 4190
rect 16960 4170 16970 4190
rect 16990 4170 17060 4190
rect 17080 4170 17090 4190
rect 17140 4170 17150 4190
rect 17170 4170 17240 4190
rect 17260 4170 17270 4190
rect 17320 4170 17330 4190
rect 17350 4170 17420 4190
rect 17440 4170 17450 4190
rect 17500 4170 17510 4190
rect 17530 4170 17600 4190
rect 17620 4170 17630 4190
rect 17680 4170 17690 4190
rect 17710 4170 17780 4190
rect 17800 4170 17810 4190
rect 17860 4170 17870 4190
rect 17890 4170 17960 4190
rect 17980 4170 17990 4190
rect 18040 4170 18050 4190
rect 18070 4170 18140 4190
rect 18160 4170 18170 4190
rect 18220 4170 18230 4190
rect 18250 4170 18320 4190
rect 18340 4170 18350 4190
rect 18400 4170 18410 4190
rect 18430 4170 18500 4190
rect 18520 4170 18530 4190
rect 18580 4170 18590 4190
rect 18610 4170 18680 4190
rect 18700 4170 18710 4190
rect 18760 4170 18770 4190
rect 18790 4170 18860 4190
rect 18880 4170 18890 4190
rect 18940 4170 18950 4190
rect 18970 4170 19040 4190
rect 19060 4170 19070 4190
rect 19120 4170 19130 4190
rect 19150 4170 19220 4190
rect 19240 4170 19250 4190
rect 19300 4170 19310 4190
rect 19330 4170 19400 4190
rect 19420 4170 19430 4190
rect 19480 4170 19490 4190
rect 19510 4170 19580 4190
rect 19600 4170 19610 4190
rect 19660 4170 19670 4190
rect 19690 4170 19760 4190
rect 19780 4170 19790 4190
rect 19840 4170 19850 4190
rect 19870 4170 19940 4190
rect 19960 4170 19970 4190
rect 20015 4170 20030 4190
rect 20050 4170 20120 4190
rect 20140 4170 20210 4190
rect 20230 4170 20300 4190
rect 20320 4170 20390 4190
rect 20410 4170 20480 4190
rect 20500 4170 20570 4190
rect 20590 4170 20660 4190
rect 20680 4170 20690 4190
rect 20765 4145 20785 4345
rect 9125 4125 9230 4145
rect 9250 4125 9320 4145
rect 9340 4125 9410 4145
rect 9430 4125 9500 4145
rect 9520 4125 9590 4145
rect 9610 4125 9680 4145
rect 9700 4125 9770 4145
rect 9790 4125 9860 4145
rect 9880 4125 9950 4145
rect 9970 4125 10040 4145
rect 10060 4125 10130 4145
rect 10150 4125 10220 4145
rect 10240 4125 10310 4145
rect 10330 4125 10400 4145
rect 10420 4125 10490 4145
rect 10510 4125 10580 4145
rect 10600 4125 10670 4145
rect 10690 4125 10760 4145
rect 10780 4125 10850 4145
rect 10870 4125 10940 4145
rect 10960 4125 11030 4145
rect 11050 4125 11120 4145
rect 11140 4125 11210 4145
rect 11230 4125 11300 4145
rect 11320 4125 11390 4145
rect 11410 4125 11480 4145
rect 11500 4125 11570 4145
rect 11590 4125 11660 4145
rect 11680 4125 11750 4145
rect 11770 4125 11840 4145
rect 11860 4125 11930 4145
rect 11950 4125 12020 4145
rect 12040 4125 12110 4145
rect 12130 4125 12200 4145
rect 12220 4125 12290 4145
rect 12310 4125 12380 4145
rect 12400 4125 12470 4145
rect 12490 4125 12560 4145
rect 12580 4125 12650 4145
rect 12670 4125 12740 4145
rect 12760 4125 12830 4145
rect 12850 4125 12920 4145
rect 12940 4125 13010 4145
rect 13030 4125 13100 4145
rect 13120 4125 13190 4145
rect 13210 4125 13280 4145
rect 13300 4125 13370 4145
rect 13390 4125 13460 4145
rect 13480 4125 13550 4145
rect 13570 4125 13640 4145
rect 13660 4125 13730 4145
rect 13750 4125 13820 4145
rect 13840 4125 13910 4145
rect 13930 4125 14000 4145
rect 14020 4125 14090 4145
rect 14110 4125 14180 4145
rect 14200 4125 14270 4145
rect 14290 4125 14360 4145
rect 14380 4125 14450 4145
rect 14470 4125 14540 4145
rect 14560 4125 14630 4145
rect 14650 4125 14720 4145
rect 14740 4125 14810 4145
rect 14830 4125 14900 4145
rect 14920 4125 14990 4145
rect 15010 4125 15080 4145
rect 15100 4125 15170 4145
rect 15190 4125 15260 4145
rect 15280 4125 15350 4145
rect 15370 4125 15440 4145
rect 15460 4125 15530 4145
rect 15550 4125 15620 4145
rect 15640 4125 15710 4145
rect 15730 4125 15800 4145
rect 15820 4125 15890 4145
rect 15910 4125 15980 4145
rect 16000 4125 16070 4145
rect 16090 4125 16160 4145
rect 16180 4125 16250 4145
rect 16270 4125 16340 4145
rect 16360 4125 16430 4145
rect 16450 4125 16520 4145
rect 16540 4125 16610 4145
rect 16630 4125 16700 4145
rect 16720 4125 16790 4145
rect 16810 4125 16880 4145
rect 16900 4125 16970 4145
rect 16990 4125 17060 4145
rect 17080 4125 17150 4145
rect 17170 4125 17240 4145
rect 17260 4125 17330 4145
rect 17350 4125 17420 4145
rect 17440 4125 17510 4145
rect 17530 4125 17600 4145
rect 17620 4125 17690 4145
rect 17710 4125 17780 4145
rect 17800 4125 17870 4145
rect 17890 4125 17960 4145
rect 17980 4125 18050 4145
rect 18070 4125 18140 4145
rect 18160 4125 18230 4145
rect 18250 4125 18320 4145
rect 18340 4125 18410 4145
rect 18430 4125 18500 4145
rect 18520 4125 18590 4145
rect 18610 4125 18680 4145
rect 18700 4125 18770 4145
rect 18790 4125 18860 4145
rect 18880 4125 18950 4145
rect 18970 4125 19040 4145
rect 19060 4125 19130 4145
rect 19150 4125 19220 4145
rect 19240 4125 19310 4145
rect 19330 4125 19400 4145
rect 19420 4125 19490 4145
rect 19510 4125 19580 4145
rect 19600 4125 19670 4145
rect 19690 4125 19760 4145
rect 19780 4125 19850 4145
rect 19870 4125 19940 4145
rect 19960 4125 20030 4145
rect 20050 4125 20120 4145
rect 20140 4125 20210 4145
rect 20230 4125 20300 4145
rect 20320 4125 20390 4145
rect 20410 4125 20480 4145
rect 20500 4125 20570 4145
rect 20590 4125 20660 4145
rect 20680 4125 20785 4145
rect 9175 4085 10040 4105
rect 10060 4085 10580 4105
rect 10600 4085 10760 4105
rect 10780 4085 11300 4105
rect 11320 4085 11480 4105
rect 11500 4085 12020 4105
rect 12040 4085 12200 4105
rect 12220 4085 12740 4105
rect 12760 4085 12920 4105
rect 12940 4085 13460 4105
rect 13480 4085 13640 4105
rect 13660 4085 13775 4105
rect 13795 4085 13865 4105
rect 13885 4085 13955 4105
rect 13975 4085 14180 4105
rect 14200 4085 15710 4105
rect 15730 4085 15935 4105
rect 15955 4085 16025 4105
rect 16045 4085 16115 4105
rect 16135 4085 16250 4105
rect 16270 4085 16430 4105
rect 16450 4085 16970 4105
rect 16990 4085 17150 4105
rect 17170 4085 17690 4105
rect 17710 4085 17870 4105
rect 17890 4085 18410 4105
rect 18430 4085 18590 4105
rect 18610 4085 19130 4105
rect 19150 4085 19310 4105
rect 19330 4085 19850 4105
rect 19870 4085 20735 4105
rect 20840 4065 20860 4375
rect 9050 4045 9230 4065
rect 9250 4045 9320 4065
rect 9340 4045 9410 4065
rect 9430 4045 9500 4065
rect 9520 4045 9590 4065
rect 9610 4045 9680 4065
rect 9700 4045 9770 4065
rect 9790 4045 9860 4065
rect 9880 4045 9950 4065
rect 9970 4045 10040 4065
rect 10060 4045 10130 4065
rect 10150 4045 10220 4065
rect 10240 4045 10310 4065
rect 10330 4045 10400 4065
rect 10420 4045 10490 4065
rect 10510 4045 10580 4065
rect 10600 4045 10670 4065
rect 10690 4045 10760 4065
rect 10780 4045 10850 4065
rect 10870 4045 10940 4065
rect 10960 4045 11030 4065
rect 11050 4045 11120 4065
rect 11140 4045 11210 4065
rect 11230 4045 11300 4065
rect 11320 4045 11390 4065
rect 11410 4045 11480 4065
rect 11500 4045 11570 4065
rect 11590 4045 11660 4065
rect 11680 4045 11750 4065
rect 11770 4045 11840 4065
rect 11860 4045 11930 4065
rect 11950 4045 12020 4065
rect 12040 4045 12110 4065
rect 12130 4045 12200 4065
rect 12220 4045 12290 4065
rect 12310 4045 12380 4065
rect 12400 4045 12470 4065
rect 12490 4045 12560 4065
rect 12580 4045 12650 4065
rect 12670 4045 12740 4065
rect 12760 4045 12830 4065
rect 12850 4045 12920 4065
rect 12940 4045 13010 4065
rect 13030 4045 13100 4065
rect 13120 4045 13190 4065
rect 13210 4045 13280 4065
rect 13300 4045 13370 4065
rect 13390 4045 13460 4065
rect 13480 4045 13550 4065
rect 13570 4045 13640 4065
rect 13660 4045 13730 4065
rect 13750 4045 13820 4065
rect 13840 4045 13910 4065
rect 13930 4045 14000 4065
rect 14020 4045 14090 4065
rect 14110 4045 14180 4065
rect 14200 4045 14270 4065
rect 14290 4045 14360 4065
rect 14380 4045 14450 4065
rect 14470 4045 14540 4065
rect 14560 4045 14630 4065
rect 14650 4045 14720 4065
rect 14740 4045 14810 4065
rect 14830 4045 14900 4065
rect 14920 4045 14990 4065
rect 15010 4045 15080 4065
rect 15100 4045 15170 4065
rect 15190 4045 15260 4065
rect 15280 4045 15350 4065
rect 15370 4045 15440 4065
rect 15460 4045 15530 4065
rect 15550 4045 15620 4065
rect 15640 4045 15710 4065
rect 15730 4045 15800 4065
rect 15820 4045 15890 4065
rect 15910 4045 15980 4065
rect 16000 4045 16070 4065
rect 16090 4045 16160 4065
rect 16180 4045 16250 4065
rect 16270 4045 16340 4065
rect 16360 4045 16430 4065
rect 16450 4045 16520 4065
rect 16540 4045 16610 4065
rect 16630 4045 16700 4065
rect 16720 4045 16790 4065
rect 16810 4045 16880 4065
rect 16900 4045 16970 4065
rect 16990 4045 17060 4065
rect 17080 4045 17150 4065
rect 17170 4045 17240 4065
rect 17260 4045 17330 4065
rect 17350 4045 17420 4065
rect 17440 4045 17510 4065
rect 17530 4045 17600 4065
rect 17620 4045 17690 4065
rect 17710 4045 17780 4065
rect 17800 4045 17870 4065
rect 17890 4045 17960 4065
rect 17980 4045 18050 4065
rect 18070 4045 18140 4065
rect 18160 4045 18230 4065
rect 18250 4045 18320 4065
rect 18340 4045 18410 4065
rect 18430 4045 18500 4065
rect 18520 4045 18590 4065
rect 18610 4045 18680 4065
rect 18700 4045 18770 4065
rect 18790 4045 18860 4065
rect 18880 4045 18950 4065
rect 18970 4045 19040 4065
rect 19060 4045 19130 4065
rect 19150 4045 19220 4065
rect 19240 4045 19310 4065
rect 19330 4045 19400 4065
rect 19420 4045 19490 4065
rect 19510 4045 19580 4065
rect 19600 4045 19670 4065
rect 19690 4045 19760 4065
rect 19780 4045 19850 4065
rect 19870 4045 19940 4065
rect 19960 4045 20030 4065
rect 20050 4045 20120 4065
rect 20140 4045 20210 4065
rect 20230 4045 20300 4065
rect 20320 4045 20390 4065
rect 20410 4045 20480 4065
rect 20500 4045 20570 4065
rect 20590 4045 20660 4065
rect 20680 4045 20860 4065
rect 9175 4005 13550 4025
rect 13570 4005 14090 4025
rect 14110 4005 15800 4025
rect 15820 4005 16340 4025
rect 16360 4005 20345 4025
rect 20365 4005 20735 4025
rect 9175 3965 13730 3985
rect 13750 3965 13910 3985
rect 13930 3965 15980 3985
rect 16000 3965 16160 3985
rect 16180 3965 20435 3985
rect 20455 3965 20735 3985
rect 9175 3925 10085 3945
rect 10105 3925 10265 3945
rect 10285 3925 10445 3945
rect 10465 3925 10805 3945
rect 10825 3925 10985 3945
rect 11005 3925 11165 3945
rect 11185 3925 11525 3945
rect 11545 3925 11705 3945
rect 11725 3925 11885 3945
rect 11905 3925 12245 3945
rect 12265 3925 12425 3945
rect 12445 3925 12605 3945
rect 12625 3925 12965 3945
rect 12985 3925 13145 3945
rect 13165 3925 13325 3945
rect 13345 3925 14405 3945
rect 14425 3925 14585 3945
rect 14605 3925 14765 3945
rect 14785 3925 15125 3945
rect 15145 3925 15305 3945
rect 15325 3925 15485 3945
rect 15505 3925 16565 3945
rect 16585 3925 16745 3945
rect 16765 3925 16925 3945
rect 16945 3925 17285 3945
rect 17305 3925 17465 3945
rect 17485 3925 17645 3945
rect 17665 3925 18005 3945
rect 18025 3925 18185 3945
rect 18205 3925 18365 3945
rect 18385 3925 18725 3945
rect 18745 3925 18905 3945
rect 18925 3925 19085 3945
rect 19105 3925 19445 3945
rect 19465 3925 19625 3945
rect 19645 3925 19805 3945
rect 19825 3925 20735 3945
rect 9175 3885 10130 3905
rect 10150 3885 10175 3905
rect 10195 3885 10220 3905
rect 10240 3885 10310 3905
rect 10330 3885 10355 3905
rect 10375 3885 10400 3905
rect 10420 3885 10850 3905
rect 10870 3885 10895 3905
rect 10915 3885 10940 3905
rect 10960 3885 11030 3905
rect 11050 3885 11075 3905
rect 11095 3885 11120 3905
rect 11140 3885 11570 3905
rect 11590 3885 11615 3905
rect 11635 3885 11660 3905
rect 11680 3885 11750 3905
rect 11770 3885 11795 3905
rect 11815 3885 11840 3905
rect 11860 3885 12290 3905
rect 12310 3885 12335 3905
rect 12355 3885 12380 3905
rect 12400 3885 12470 3905
rect 12490 3885 12515 3905
rect 12535 3885 12560 3905
rect 12580 3885 13010 3905
rect 13030 3885 13055 3905
rect 13075 3885 13100 3905
rect 13120 3885 13190 3905
rect 13210 3885 13235 3905
rect 13255 3885 13280 3905
rect 13300 3885 16610 3905
rect 16630 3885 16655 3905
rect 16675 3885 16700 3905
rect 16720 3885 16790 3905
rect 16810 3885 16835 3905
rect 16855 3885 16880 3905
rect 16900 3885 17330 3905
rect 17350 3885 17375 3905
rect 17395 3885 17420 3905
rect 17440 3885 17510 3905
rect 17530 3885 17555 3905
rect 17575 3885 17600 3905
rect 17620 3885 18050 3905
rect 18070 3885 18095 3905
rect 18115 3885 18140 3905
rect 18160 3885 18230 3905
rect 18250 3885 18275 3905
rect 18295 3885 18320 3905
rect 18340 3885 18770 3905
rect 18790 3885 18815 3905
rect 18835 3885 18860 3905
rect 18880 3885 18950 3905
rect 18970 3885 18995 3905
rect 19015 3885 19040 3905
rect 19060 3885 19490 3905
rect 19510 3885 19535 3905
rect 19555 3885 19580 3905
rect 19600 3885 19670 3905
rect 19690 3885 19715 3905
rect 19735 3885 19760 3905
rect 19780 3885 20735 3905
rect 9175 3845 13820 3865
rect 13840 3845 14000 3865
rect 14020 3845 14450 3865
rect 14470 3845 14630 3865
rect 14650 3845 15260 3865
rect 15280 3845 15440 3865
rect 15460 3845 15890 3865
rect 15910 3845 16070 3865
rect 16090 3845 20735 3865
rect 9175 3805 10085 3825
rect 10105 3805 10265 3825
rect 10285 3805 10445 3825
rect 10465 3805 10805 3825
rect 10825 3805 10985 3825
rect 11005 3805 11165 3825
rect 11185 3805 11525 3825
rect 11545 3805 11705 3825
rect 11725 3805 11885 3825
rect 11905 3805 12245 3825
rect 12265 3805 12425 3825
rect 12445 3805 12605 3825
rect 12625 3805 12965 3825
rect 12985 3805 13145 3825
rect 13165 3805 13325 3825
rect 13345 3805 13685 3825
rect 13705 3805 13865 3825
rect 13885 3805 14045 3825
rect 14065 3805 15845 3825
rect 15865 3805 16025 3825
rect 16045 3805 16205 3825
rect 16225 3805 16565 3825
rect 16585 3805 16745 3825
rect 16765 3805 16925 3825
rect 16945 3805 17285 3825
rect 17305 3805 17465 3825
rect 17485 3805 17645 3825
rect 17665 3805 18005 3825
rect 18025 3805 18185 3825
rect 18205 3805 18365 3825
rect 18385 3805 18725 3825
rect 18745 3805 18905 3825
rect 18925 3805 19085 3825
rect 19105 3805 19445 3825
rect 19465 3805 19625 3825
rect 19645 3805 19805 3825
rect 19825 3805 20735 3825
rect 9175 3765 9950 3785
rect 9970 3765 10490 3785
rect 10510 3765 10670 3785
rect 10690 3765 11210 3785
rect 11230 3765 11390 3785
rect 11410 3765 11930 3785
rect 11950 3765 12110 3785
rect 12130 3765 12650 3785
rect 12670 3765 12830 3785
rect 12850 3765 13370 3785
rect 13390 3765 14270 3785
rect 14290 3765 14495 3785
rect 14515 3765 14585 3785
rect 14605 3765 14675 3785
rect 14695 3765 14810 3785
rect 14830 3765 15080 3785
rect 15100 3765 15215 3785
rect 15235 3765 15305 3785
rect 15325 3765 15395 3785
rect 15415 3765 15620 3785
rect 15640 3765 16520 3785
rect 16540 3765 17060 3785
rect 17080 3765 17240 3785
rect 17260 3765 17780 3785
rect 17800 3765 17960 3785
rect 17980 3765 18500 3785
rect 18520 3765 18680 3785
rect 18700 3765 19220 3785
rect 19240 3765 19400 3785
rect 19420 3765 19940 3785
rect 19960 3765 20735 3785
rect 9175 3725 14540 3745
rect 14560 3725 14720 3745
rect 14740 3725 15170 3745
rect 15190 3725 15350 3745
rect 15370 3725 20615 3745
rect 20635 3725 20735 3745
rect 9175 3685 14360 3705
rect 14380 3685 14900 3705
rect 14920 3685 14990 3705
rect 15010 3685 15530 3705
rect 15550 3685 20525 3705
rect 20545 3685 20735 3705
rect 9050 3645 9230 3665
rect 9250 3645 9320 3665
rect 9340 3645 9410 3665
rect 9430 3645 9500 3665
rect 9520 3645 9590 3665
rect 9610 3645 9680 3665
rect 9700 3645 9770 3665
rect 9790 3645 9860 3665
rect 9880 3645 9950 3665
rect 9970 3645 10040 3665
rect 10060 3645 10130 3665
rect 10150 3645 10220 3665
rect 10240 3645 10310 3665
rect 10330 3645 10400 3665
rect 10420 3645 10490 3665
rect 10510 3645 10580 3665
rect 10600 3645 10670 3665
rect 10690 3645 10760 3665
rect 10780 3645 10850 3665
rect 10870 3645 10940 3665
rect 10960 3645 11030 3665
rect 11050 3645 11120 3665
rect 11140 3645 11210 3665
rect 11230 3645 11300 3665
rect 11320 3645 11390 3665
rect 11410 3645 11480 3665
rect 11500 3645 11570 3665
rect 11590 3645 11660 3665
rect 11680 3645 11750 3665
rect 11770 3645 11840 3665
rect 11860 3645 11930 3665
rect 11950 3645 12020 3665
rect 12040 3645 12110 3665
rect 12130 3645 12200 3665
rect 12220 3645 12290 3665
rect 12310 3645 12380 3665
rect 12400 3645 12470 3665
rect 12490 3645 12560 3665
rect 12580 3645 12650 3665
rect 12670 3645 12740 3665
rect 12760 3645 12830 3665
rect 12850 3645 12920 3665
rect 12940 3645 13010 3665
rect 13030 3645 13100 3665
rect 13120 3645 13190 3665
rect 13210 3645 13280 3665
rect 13300 3645 13370 3665
rect 13390 3645 13460 3665
rect 13480 3645 13550 3665
rect 13570 3645 13640 3665
rect 13660 3645 13730 3665
rect 13750 3645 13820 3665
rect 13840 3645 13910 3665
rect 13930 3645 14000 3665
rect 14020 3645 14090 3665
rect 14110 3645 14180 3665
rect 14200 3645 14270 3665
rect 14290 3645 14360 3665
rect 14380 3645 14450 3665
rect 14470 3645 14540 3665
rect 14560 3645 14630 3665
rect 14650 3645 14720 3665
rect 14740 3645 14810 3665
rect 14830 3645 14900 3665
rect 14920 3645 14990 3665
rect 15010 3645 15080 3665
rect 15100 3645 15170 3665
rect 15190 3645 15260 3665
rect 15280 3645 15350 3665
rect 15370 3645 15440 3665
rect 15460 3645 15530 3665
rect 15550 3645 15620 3665
rect 15640 3645 15710 3665
rect 15730 3645 15800 3665
rect 15820 3645 15890 3665
rect 15910 3645 15980 3665
rect 16000 3645 16070 3665
rect 16090 3645 16160 3665
rect 16180 3645 16250 3665
rect 16270 3645 16340 3665
rect 16360 3645 16430 3665
rect 16450 3645 16520 3665
rect 16540 3645 16610 3665
rect 16630 3645 16700 3665
rect 16720 3645 16790 3665
rect 16810 3645 16880 3665
rect 16900 3645 16970 3665
rect 16990 3645 17060 3665
rect 17080 3645 17150 3665
rect 17170 3645 17240 3665
rect 17260 3645 17330 3665
rect 17350 3645 17420 3665
rect 17440 3645 17510 3665
rect 17530 3645 17600 3665
rect 17620 3645 17690 3665
rect 17710 3645 17780 3665
rect 17800 3645 17870 3665
rect 17890 3645 17960 3665
rect 17980 3645 18050 3665
rect 18070 3645 18140 3665
rect 18160 3645 18230 3665
rect 18250 3645 18320 3665
rect 18340 3645 18410 3665
rect 18430 3645 18500 3665
rect 18520 3645 18590 3665
rect 18610 3645 18680 3665
rect 18700 3645 18770 3665
rect 18790 3645 18860 3665
rect 18880 3645 18950 3665
rect 18970 3645 19040 3665
rect 19060 3645 19130 3665
rect 19150 3645 19220 3665
rect 19240 3645 19310 3665
rect 19330 3645 19400 3665
rect 19420 3645 19490 3665
rect 19510 3645 19580 3665
rect 19600 3645 19670 3665
rect 19690 3645 19760 3665
rect 19780 3645 19850 3665
rect 19870 3645 19940 3665
rect 19960 3645 20030 3665
rect 20050 3645 20120 3665
rect 20140 3645 20210 3665
rect 20230 3645 20300 3665
rect 20320 3645 20390 3665
rect 20410 3645 20480 3665
rect 20500 3645 20570 3665
rect 20590 3645 20660 3665
rect 20680 3645 20860 3665
rect 9050 3445 9070 3645
rect 9220 3600 9230 3620
rect 9250 3600 9320 3620
rect 9340 3600 9410 3620
rect 9430 3600 9500 3620
rect 9520 3600 9590 3620
rect 9610 3600 9680 3620
rect 9700 3600 9770 3620
rect 9790 3600 9860 3620
rect 9880 3600 9890 3620
rect 9940 3600 9950 3620
rect 9970 3600 10040 3620
rect 10060 3600 10070 3620
rect 10120 3600 10130 3620
rect 10150 3600 10220 3620
rect 10240 3600 10250 3620
rect 10300 3600 10310 3620
rect 10330 3600 10400 3620
rect 10420 3600 10430 3620
rect 10480 3600 10490 3620
rect 10510 3600 10580 3620
rect 10600 3600 10610 3620
rect 10660 3600 10670 3620
rect 10690 3600 10760 3620
rect 10780 3600 10790 3620
rect 10840 3600 10850 3620
rect 10870 3600 10940 3620
rect 10960 3600 10970 3620
rect 11020 3600 11030 3620
rect 11050 3600 11120 3620
rect 11140 3600 11150 3620
rect 11200 3600 11210 3620
rect 11230 3600 11300 3620
rect 11320 3600 11330 3620
rect 11380 3600 11390 3620
rect 11410 3600 11480 3620
rect 11500 3600 11510 3620
rect 11560 3600 11570 3620
rect 11590 3600 11660 3620
rect 11680 3600 11690 3620
rect 11740 3600 11750 3620
rect 11770 3600 11840 3620
rect 11860 3600 11870 3620
rect 11920 3600 11930 3620
rect 11950 3600 12020 3620
rect 12040 3600 12050 3620
rect 12100 3600 12110 3620
rect 12130 3600 12200 3620
rect 12220 3600 12230 3620
rect 12280 3600 12290 3620
rect 12310 3600 12380 3620
rect 12400 3600 12410 3620
rect 12460 3600 12470 3620
rect 12490 3600 12560 3620
rect 12580 3600 12590 3620
rect 12640 3600 12650 3620
rect 12670 3600 12740 3620
rect 12760 3600 12770 3620
rect 12820 3600 12830 3620
rect 12850 3600 12920 3620
rect 12940 3600 12950 3620
rect 13000 3600 13010 3620
rect 13030 3600 13100 3620
rect 13120 3600 13130 3620
rect 13180 3600 13190 3620
rect 13210 3600 13280 3620
rect 13300 3600 13310 3620
rect 13360 3600 13370 3620
rect 13390 3600 13460 3620
rect 13480 3600 13490 3620
rect 13540 3600 13550 3620
rect 13570 3600 13640 3620
rect 13660 3600 13670 3620
rect 13720 3600 13730 3620
rect 13750 3600 13820 3620
rect 13840 3600 13850 3620
rect 13900 3600 13910 3620
rect 13930 3600 14000 3620
rect 14020 3600 14030 3620
rect 14080 3600 14090 3620
rect 14110 3600 14180 3620
rect 14200 3600 14210 3620
rect 14260 3600 14270 3620
rect 14290 3600 14360 3620
rect 14380 3600 14390 3620
rect 14440 3600 14450 3620
rect 14470 3600 14540 3620
rect 14560 3600 14570 3620
rect 14620 3600 14630 3620
rect 14650 3600 14720 3620
rect 14740 3600 14750 3620
rect 14800 3600 14810 3620
rect 14830 3600 14900 3620
rect 14920 3600 14930 3620
rect 14980 3600 14990 3620
rect 15010 3600 15080 3620
rect 15100 3600 15110 3620
rect 15160 3600 15170 3620
rect 15190 3600 15260 3620
rect 15280 3600 15290 3620
rect 15340 3600 15350 3620
rect 15370 3600 15440 3620
rect 15460 3600 15470 3620
rect 15520 3600 15530 3620
rect 15550 3600 15620 3620
rect 15640 3600 15650 3620
rect 15700 3600 15710 3620
rect 15730 3600 15800 3620
rect 15820 3600 15830 3620
rect 15880 3600 15890 3620
rect 15910 3600 15980 3620
rect 16000 3600 16010 3620
rect 16060 3600 16070 3620
rect 16090 3600 16160 3620
rect 16180 3600 16190 3620
rect 16240 3600 16250 3620
rect 16270 3600 16340 3620
rect 16360 3600 16370 3620
rect 16420 3600 16430 3620
rect 16450 3600 16520 3620
rect 16540 3600 16550 3620
rect 16600 3600 16610 3620
rect 16630 3600 16700 3620
rect 16720 3600 16730 3620
rect 16780 3600 16790 3620
rect 16810 3600 16880 3620
rect 16900 3600 16910 3620
rect 16960 3600 16970 3620
rect 16990 3600 17060 3620
rect 17080 3600 17090 3620
rect 17140 3600 17150 3620
rect 17170 3600 17240 3620
rect 17260 3600 17270 3620
rect 17320 3600 17330 3620
rect 17350 3600 17420 3620
rect 17440 3600 17450 3620
rect 17500 3600 17510 3620
rect 17530 3600 17600 3620
rect 17620 3600 17630 3620
rect 17680 3600 17690 3620
rect 17710 3600 17780 3620
rect 17800 3600 17810 3620
rect 17860 3600 17870 3620
rect 17890 3600 17960 3620
rect 17980 3600 17990 3620
rect 18040 3600 18050 3620
rect 18070 3600 18140 3620
rect 18160 3600 18170 3620
rect 18220 3600 18230 3620
rect 18250 3600 18320 3620
rect 18340 3600 18350 3620
rect 18400 3600 18410 3620
rect 18430 3600 18500 3620
rect 18520 3600 18530 3620
rect 18580 3600 18590 3620
rect 18610 3600 18680 3620
rect 18700 3600 18710 3620
rect 18760 3600 18770 3620
rect 18790 3600 18860 3620
rect 18880 3600 18890 3620
rect 18940 3600 18950 3620
rect 18970 3600 19040 3620
rect 19060 3600 19070 3620
rect 19120 3600 19130 3620
rect 19150 3600 19220 3620
rect 19240 3600 19250 3620
rect 19300 3600 19310 3620
rect 19330 3600 19400 3620
rect 19420 3600 19430 3620
rect 19480 3600 19490 3620
rect 19510 3600 19580 3620
rect 19600 3600 19610 3620
rect 19660 3600 19670 3620
rect 19690 3600 19760 3620
rect 19780 3600 19790 3620
rect 19840 3600 19850 3620
rect 19870 3600 19940 3620
rect 19960 3600 19970 3620
rect 20020 3600 20030 3620
rect 20050 3600 20120 3620
rect 20140 3600 20210 3620
rect 20230 3600 20300 3620
rect 20320 3600 20390 3620
rect 20410 3600 20480 3620
rect 20500 3600 20570 3620
rect 20590 3600 20660 3620
rect 20680 3600 20690 3620
rect 9185 3565 9205 3575
rect 9185 3475 9205 3485
rect 9275 3565 9295 3575
rect 9275 3475 9295 3485
rect 9365 3565 9385 3575
rect 9365 3475 9385 3485
rect 9455 3565 9475 3600
rect 9455 3475 9475 3485
rect 9545 3565 9565 3575
rect 9545 3475 9565 3485
rect 9635 3565 9655 3600
rect 9635 3475 9655 3485
rect 9725 3565 9745 3575
rect 9725 3475 9745 3485
rect 9815 3565 9835 3575
rect 9815 3475 9835 3485
rect 9905 3565 9925 3575
rect 9905 3475 9925 3485
rect 9995 3565 10015 3575
rect 9995 3475 10015 3485
rect 10085 3565 10105 3575
rect 10085 3475 10105 3485
rect 10175 3565 10195 3575
rect 10175 3475 10195 3485
rect 10265 3565 10285 3575
rect 10265 3475 10285 3485
rect 10355 3565 10375 3575
rect 10355 3475 10375 3485
rect 10445 3565 10465 3575
rect 10445 3475 10465 3485
rect 10535 3565 10555 3575
rect 10535 3475 10555 3485
rect 10625 3565 10645 3575
rect 10625 3475 10645 3485
rect 10715 3565 10735 3575
rect 10715 3475 10735 3485
rect 10805 3565 10825 3575
rect 10805 3475 10825 3485
rect 10895 3565 10915 3575
rect 10895 3475 10915 3485
rect 10985 3565 11005 3575
rect 10985 3475 11005 3485
rect 11075 3565 11095 3575
rect 11075 3475 11095 3485
rect 11165 3565 11185 3575
rect 11165 3475 11185 3485
rect 11255 3565 11275 3575
rect 11255 3475 11275 3485
rect 11345 3565 11365 3575
rect 11345 3475 11365 3485
rect 11435 3565 11455 3575
rect 11435 3475 11455 3485
rect 11525 3565 11545 3575
rect 11525 3475 11545 3485
rect 11615 3565 11635 3575
rect 11615 3475 11635 3485
rect 11705 3565 11725 3575
rect 11705 3475 11725 3485
rect 11795 3565 11815 3575
rect 11795 3475 11815 3485
rect 11885 3565 11905 3575
rect 11885 3475 11905 3485
rect 11975 3565 11995 3575
rect 11975 3475 11995 3485
rect 12065 3565 12085 3575
rect 12065 3475 12085 3485
rect 12155 3565 12175 3575
rect 12155 3475 12175 3485
rect 12245 3565 12265 3575
rect 12245 3475 12265 3485
rect 12335 3565 12355 3575
rect 12335 3475 12355 3485
rect 12425 3565 12445 3575
rect 12425 3475 12445 3485
rect 12515 3565 12535 3575
rect 12515 3475 12535 3485
rect 12605 3565 12625 3575
rect 12605 3475 12625 3485
rect 12695 3565 12715 3575
rect 12695 3475 12715 3485
rect 12785 3565 12805 3575
rect 12785 3475 12805 3485
rect 12875 3565 12895 3575
rect 12875 3475 12895 3485
rect 12965 3565 12985 3575
rect 12965 3475 12985 3485
rect 13055 3565 13075 3575
rect 13055 3475 13075 3485
rect 13145 3565 13165 3575
rect 13145 3475 13165 3485
rect 13235 3565 13255 3575
rect 13235 3475 13255 3485
rect 13325 3565 13345 3575
rect 13325 3475 13345 3485
rect 13415 3565 13435 3575
rect 13415 3475 13435 3485
rect 13505 3565 13525 3575
rect 13505 3475 13525 3485
rect 13595 3565 13615 3575
rect 13595 3475 13615 3485
rect 13685 3565 13705 3575
rect 13685 3475 13705 3485
rect 13775 3565 13795 3575
rect 13775 3475 13795 3485
rect 13865 3565 13885 3575
rect 13865 3475 13885 3485
rect 13955 3565 13975 3575
rect 13955 3475 13975 3485
rect 14045 3565 14065 3575
rect 14045 3475 14065 3485
rect 14135 3565 14155 3575
rect 14135 3475 14155 3485
rect 14225 3565 14245 3575
rect 14225 3475 14245 3485
rect 14315 3565 14335 3575
rect 14315 3475 14335 3485
rect 14405 3565 14425 3575
rect 14405 3475 14425 3485
rect 14495 3565 14515 3575
rect 14495 3475 14515 3485
rect 14585 3565 14605 3575
rect 14585 3475 14605 3485
rect 14675 3565 14695 3575
rect 14675 3475 14695 3485
rect 14765 3565 14785 3575
rect 14765 3475 14785 3485
rect 14855 3565 14875 3575
rect 14855 3475 14875 3485
rect 14945 3565 14965 3575
rect 14945 3475 14965 3485
rect 15035 3565 15055 3575
rect 15035 3475 15055 3485
rect 15125 3565 15145 3575
rect 15125 3475 15145 3485
rect 15215 3565 15235 3575
rect 15215 3475 15235 3485
rect 15305 3565 15325 3575
rect 15305 3475 15325 3485
rect 15395 3565 15415 3575
rect 15395 3475 15415 3485
rect 15485 3565 15505 3575
rect 15485 3475 15505 3485
rect 15575 3565 15595 3575
rect 15575 3475 15595 3485
rect 15665 3565 15685 3575
rect 15665 3475 15685 3485
rect 15755 3565 15775 3575
rect 15755 3475 15775 3485
rect 15845 3565 15865 3575
rect 15845 3475 15865 3485
rect 15935 3565 15955 3575
rect 15935 3475 15955 3485
rect 16025 3565 16045 3575
rect 16025 3475 16045 3485
rect 16115 3565 16135 3575
rect 16115 3475 16135 3485
rect 16205 3565 16225 3575
rect 16205 3475 16225 3485
rect 16295 3565 16315 3575
rect 16295 3475 16315 3485
rect 16385 3565 16405 3575
rect 16385 3475 16405 3485
rect 16475 3565 16495 3575
rect 16475 3475 16495 3485
rect 16565 3565 16585 3575
rect 16565 3475 16585 3485
rect 16655 3565 16675 3575
rect 16655 3475 16675 3485
rect 16745 3565 16765 3575
rect 16745 3475 16765 3485
rect 16835 3565 16855 3575
rect 16835 3475 16855 3485
rect 16925 3565 16945 3575
rect 16925 3475 16945 3485
rect 17015 3565 17035 3575
rect 17015 3475 17035 3485
rect 17105 3565 17125 3575
rect 17105 3475 17125 3485
rect 17195 3565 17215 3575
rect 17195 3475 17215 3485
rect 17285 3565 17305 3575
rect 17285 3475 17305 3485
rect 17375 3565 17395 3575
rect 17375 3475 17395 3485
rect 17465 3565 17485 3575
rect 17465 3475 17485 3485
rect 17555 3565 17575 3575
rect 17555 3475 17575 3485
rect 17645 3565 17665 3575
rect 17645 3475 17665 3485
rect 17735 3565 17755 3575
rect 17735 3475 17755 3485
rect 17825 3565 17845 3575
rect 17825 3475 17845 3485
rect 17915 3565 17935 3575
rect 17915 3475 17935 3485
rect 18005 3565 18025 3575
rect 18005 3475 18025 3485
rect 18095 3565 18115 3575
rect 18095 3475 18115 3485
rect 18185 3565 18205 3575
rect 18185 3475 18205 3485
rect 18275 3565 18295 3575
rect 18275 3475 18295 3485
rect 18365 3565 18385 3575
rect 18365 3475 18385 3485
rect 18455 3565 18475 3575
rect 18455 3475 18475 3485
rect 18545 3565 18565 3575
rect 18545 3475 18565 3485
rect 18635 3565 18655 3575
rect 18635 3475 18655 3485
rect 18725 3565 18745 3575
rect 18725 3475 18745 3485
rect 18815 3565 18835 3575
rect 18815 3475 18835 3485
rect 18905 3565 18925 3575
rect 18905 3475 18925 3485
rect 18995 3565 19015 3575
rect 18995 3475 19015 3485
rect 19085 3565 19105 3575
rect 19085 3475 19105 3485
rect 19175 3565 19195 3575
rect 19175 3475 19195 3485
rect 19265 3565 19285 3575
rect 19265 3475 19285 3485
rect 19355 3565 19375 3575
rect 19355 3475 19375 3485
rect 19445 3565 19465 3575
rect 19445 3475 19465 3485
rect 19535 3565 19555 3575
rect 19535 3475 19555 3485
rect 19625 3565 19645 3575
rect 19625 3475 19645 3485
rect 19715 3565 19735 3575
rect 19715 3475 19735 3485
rect 19805 3565 19825 3575
rect 19805 3475 19825 3485
rect 19895 3565 19915 3575
rect 19895 3475 19915 3485
rect 19985 3565 20005 3575
rect 19985 3475 20005 3485
rect 20075 3565 20095 3575
rect 20075 3475 20095 3485
rect 20165 3565 20185 3575
rect 20165 3475 20185 3485
rect 20255 3565 20275 3600
rect 20255 3475 20275 3485
rect 20345 3565 20365 3575
rect 20345 3475 20365 3485
rect 20435 3565 20455 3600
rect 20435 3475 20455 3485
rect 20525 3565 20545 3575
rect 20525 3475 20545 3485
rect 20615 3565 20635 3575
rect 20615 3475 20635 3485
rect 20705 3565 20725 3575
rect 20705 3475 20725 3485
rect 20840 3445 20860 3645
rect 9040 3425 9050 3445
rect 9070 3425 9185 3445
rect 9205 3425 9230 3445
rect 9250 3425 9320 3445
rect 9340 3425 9410 3445
rect 9430 3425 9500 3445
rect 9520 3425 9590 3445
rect 9610 3425 9680 3445
rect 9700 3425 9770 3445
rect 9790 3425 9860 3445
rect 9880 3425 9905 3445
rect 9925 3425 9950 3445
rect 9970 3425 10040 3445
rect 10060 3425 10085 3445
rect 10105 3425 10130 3445
rect 10150 3425 10220 3445
rect 10240 3425 10265 3445
rect 10285 3425 10310 3445
rect 10330 3425 10400 3445
rect 10420 3425 10445 3445
rect 10465 3425 10490 3445
rect 10510 3425 10580 3445
rect 10600 3425 10625 3445
rect 10645 3425 10670 3445
rect 10690 3425 10760 3445
rect 10780 3425 10805 3445
rect 10825 3425 10850 3445
rect 10870 3425 10940 3445
rect 10960 3425 10985 3445
rect 11005 3425 11030 3445
rect 11050 3425 11120 3445
rect 11140 3425 11165 3445
rect 11185 3425 11210 3445
rect 11230 3425 11300 3445
rect 11320 3425 11345 3445
rect 11365 3425 11390 3445
rect 11410 3425 11480 3445
rect 11500 3425 11525 3445
rect 11545 3425 11570 3445
rect 11590 3425 11660 3445
rect 11680 3425 11705 3445
rect 11725 3425 11750 3445
rect 11770 3425 11840 3445
rect 11860 3425 11885 3445
rect 11905 3425 11930 3445
rect 11950 3425 12020 3445
rect 12040 3425 12065 3445
rect 12085 3425 12110 3445
rect 12130 3425 12200 3445
rect 12220 3425 12245 3445
rect 12265 3425 12290 3445
rect 12310 3425 12380 3445
rect 12400 3425 12425 3445
rect 12445 3425 12470 3445
rect 12490 3425 12560 3445
rect 12580 3425 12605 3445
rect 12625 3425 12650 3445
rect 12670 3425 12740 3445
rect 12760 3425 12785 3445
rect 12805 3425 12830 3445
rect 12850 3425 12920 3445
rect 12940 3425 12965 3445
rect 12985 3425 13010 3445
rect 13030 3425 13100 3445
rect 13120 3425 13145 3445
rect 13165 3425 13190 3445
rect 13210 3425 13280 3445
rect 13300 3425 13325 3445
rect 13345 3425 13370 3445
rect 13390 3425 13460 3445
rect 13480 3425 13505 3445
rect 13525 3425 13550 3445
rect 13570 3425 13640 3445
rect 13660 3425 13685 3445
rect 13705 3425 13730 3445
rect 13750 3425 13820 3445
rect 13840 3425 13865 3445
rect 13885 3425 13910 3445
rect 13930 3425 14000 3445
rect 14020 3425 14045 3445
rect 14065 3425 14090 3445
rect 14110 3425 14180 3445
rect 14200 3425 14225 3445
rect 14245 3425 14270 3445
rect 14290 3425 14360 3445
rect 14380 3425 14405 3445
rect 14425 3425 14450 3445
rect 14470 3425 14540 3445
rect 14560 3425 14585 3445
rect 14605 3425 14630 3445
rect 14650 3425 14720 3445
rect 14740 3425 14765 3445
rect 14785 3425 14810 3445
rect 14830 3425 14900 3445
rect 14920 3425 14945 3445
rect 14965 3425 14990 3445
rect 15010 3425 15080 3445
rect 15100 3425 15125 3445
rect 15145 3425 15170 3445
rect 15190 3425 15260 3445
rect 15280 3425 15305 3445
rect 15325 3425 15350 3445
rect 15370 3425 15440 3445
rect 15460 3425 15485 3445
rect 15505 3425 15530 3445
rect 15550 3425 15620 3445
rect 15640 3425 15665 3445
rect 15685 3425 15710 3445
rect 15730 3425 15800 3445
rect 15820 3425 15845 3445
rect 15865 3425 15890 3445
rect 15910 3425 15980 3445
rect 16000 3425 16025 3445
rect 16045 3425 16070 3445
rect 16090 3425 16160 3445
rect 16180 3425 16205 3445
rect 16225 3425 16250 3445
rect 16270 3425 16340 3445
rect 16360 3425 16385 3445
rect 16405 3425 16430 3445
rect 16450 3425 16520 3445
rect 16540 3425 16565 3445
rect 16585 3425 16610 3445
rect 16630 3425 16700 3445
rect 16720 3425 16745 3445
rect 16765 3425 16790 3445
rect 16810 3425 16880 3445
rect 16900 3425 16925 3445
rect 16945 3425 16970 3445
rect 16990 3425 17060 3445
rect 17080 3425 17105 3445
rect 17125 3425 17150 3445
rect 17170 3425 17240 3445
rect 17260 3425 17285 3445
rect 17305 3425 17330 3445
rect 17350 3425 17420 3445
rect 17440 3425 17465 3445
rect 17485 3425 17510 3445
rect 17530 3425 17600 3445
rect 17620 3425 17645 3445
rect 17665 3425 17690 3445
rect 17710 3425 17780 3445
rect 17800 3425 17825 3445
rect 17845 3425 17870 3445
rect 17890 3425 17960 3445
rect 17980 3425 18005 3445
rect 18025 3425 18050 3445
rect 18070 3425 18140 3445
rect 18160 3425 18185 3445
rect 18205 3425 18230 3445
rect 18250 3425 18320 3445
rect 18340 3425 18365 3445
rect 18385 3425 18410 3445
rect 18430 3425 18500 3445
rect 18520 3425 18545 3445
rect 18565 3425 18590 3445
rect 18610 3425 18680 3445
rect 18700 3425 18725 3445
rect 18745 3425 18770 3445
rect 18790 3425 18860 3445
rect 18880 3425 18905 3445
rect 18925 3425 18950 3445
rect 18970 3425 19040 3445
rect 19060 3425 19085 3445
rect 19105 3425 19130 3445
rect 19150 3425 19220 3445
rect 19240 3425 19265 3445
rect 19285 3425 19310 3445
rect 19330 3425 19400 3445
rect 19420 3425 19445 3445
rect 19465 3425 19490 3445
rect 19510 3425 19580 3445
rect 19600 3425 19625 3445
rect 19645 3425 19670 3445
rect 19690 3425 19760 3445
rect 19780 3425 19805 3445
rect 19825 3425 19850 3445
rect 19870 3425 19940 3445
rect 19960 3425 19985 3445
rect 20005 3425 20030 3445
rect 20050 3425 20120 3445
rect 20140 3425 20210 3445
rect 20230 3425 20300 3445
rect 20320 3425 20390 3445
rect 20410 3425 20480 3445
rect 20500 3425 20570 3445
rect 20590 3425 20660 3445
rect 20680 3425 20705 3445
rect 20725 3425 20840 3445
rect 20860 3425 20870 3445
<< viali >>
rect 9185 4345 9205 4365
rect 9905 4345 9925 4365
rect 10085 4345 10105 4365
rect 10265 4345 10285 4365
rect 10445 4345 10465 4365
rect 10625 4345 10645 4365
rect 10805 4345 10825 4365
rect 10985 4345 11005 4365
rect 11165 4345 11185 4365
rect 11345 4345 11365 4365
rect 11525 4345 11545 4365
rect 11705 4345 11725 4365
rect 11885 4345 11905 4365
rect 12065 4345 12085 4365
rect 12245 4345 12265 4365
rect 12425 4345 12445 4365
rect 12605 4345 12625 4365
rect 12785 4345 12805 4365
rect 12965 4345 12985 4365
rect 13145 4345 13165 4365
rect 13325 4345 13345 4365
rect 13505 4345 13525 4365
rect 13685 4345 13705 4365
rect 13865 4345 13885 4365
rect 14045 4345 14065 4365
rect 14225 4345 14245 4365
rect 14405 4345 14425 4365
rect 14585 4345 14605 4365
rect 14765 4345 14785 4365
rect 14945 4345 14965 4365
rect 15125 4345 15145 4365
rect 15305 4345 15325 4365
rect 15485 4345 15505 4365
rect 15665 4345 15685 4365
rect 15845 4345 15865 4365
rect 16025 4345 16045 4365
rect 16205 4345 16225 4365
rect 16385 4345 16405 4365
rect 16565 4345 16585 4365
rect 16745 4345 16765 4365
rect 16925 4345 16945 4365
rect 17105 4345 17125 4365
rect 17285 4345 17305 4365
rect 17465 4345 17485 4365
rect 17645 4345 17665 4365
rect 17825 4345 17845 4365
rect 18005 4345 18025 4365
rect 18185 4345 18205 4365
rect 18365 4345 18385 4365
rect 18545 4345 18565 4365
rect 18725 4345 18745 4365
rect 18905 4345 18925 4365
rect 19085 4345 19105 4365
rect 19265 4345 19285 4365
rect 19445 4345 19465 4365
rect 19625 4345 19645 4365
rect 19805 4345 19825 4365
rect 19985 4345 20005 4365
rect 20705 4345 20725 4365
rect 9185 4225 9205 4305
rect 9905 4225 9925 4305
rect 9995 4225 10015 4305
rect 10085 4225 10105 4305
rect 10175 4225 10195 4305
rect 10265 4225 10285 4305
rect 10355 4225 10375 4305
rect 10445 4225 10465 4305
rect 10535 4225 10555 4305
rect 10625 4225 10645 4305
rect 10715 4225 10735 4305
rect 10805 4225 10825 4305
rect 10895 4225 10915 4305
rect 10985 4225 11005 4305
rect 11075 4225 11095 4305
rect 11165 4225 11185 4305
rect 11255 4225 11275 4305
rect 11345 4225 11365 4305
rect 11435 4225 11455 4305
rect 11525 4225 11545 4305
rect 11615 4225 11635 4305
rect 11705 4225 11725 4305
rect 11795 4225 11815 4305
rect 11885 4225 11905 4305
rect 11975 4225 11995 4305
rect 12065 4225 12085 4305
rect 12155 4225 12175 4305
rect 12245 4225 12265 4305
rect 12335 4225 12355 4305
rect 12425 4225 12445 4305
rect 12515 4225 12535 4305
rect 12605 4225 12625 4305
rect 12695 4225 12715 4305
rect 12785 4225 12805 4305
rect 12875 4225 12895 4305
rect 12965 4225 12985 4305
rect 13055 4225 13075 4305
rect 13145 4225 13165 4305
rect 13235 4225 13255 4305
rect 13325 4225 13345 4305
rect 13415 4225 13435 4305
rect 13505 4225 13525 4305
rect 13595 4225 13615 4305
rect 13685 4225 13705 4305
rect 13775 4225 13795 4305
rect 13865 4225 13885 4305
rect 13955 4225 13975 4305
rect 14045 4225 14065 4305
rect 14135 4225 14155 4305
rect 14225 4225 14245 4305
rect 14315 4225 14335 4305
rect 14405 4225 14425 4305
rect 14495 4225 14515 4305
rect 14585 4225 14605 4305
rect 14675 4225 14695 4305
rect 14765 4225 14785 4305
rect 14855 4225 14875 4305
rect 14945 4225 14965 4305
rect 15035 4225 15055 4305
rect 15125 4225 15145 4305
rect 15215 4225 15235 4305
rect 15305 4225 15325 4305
rect 15395 4225 15415 4305
rect 15485 4225 15505 4305
rect 15575 4225 15595 4305
rect 15665 4225 15685 4305
rect 15755 4225 15775 4305
rect 15845 4225 15865 4305
rect 15935 4225 15955 4305
rect 16025 4225 16045 4305
rect 16115 4225 16135 4305
rect 16205 4225 16225 4305
rect 16295 4225 16315 4305
rect 16385 4225 16405 4305
rect 16475 4225 16495 4305
rect 16565 4225 16585 4305
rect 16655 4225 16675 4305
rect 16745 4225 16765 4305
rect 16835 4225 16855 4305
rect 16925 4225 16945 4305
rect 17015 4225 17035 4305
rect 17105 4225 17125 4305
rect 17195 4225 17215 4305
rect 17285 4225 17305 4305
rect 17375 4225 17395 4305
rect 17465 4225 17485 4305
rect 17555 4225 17575 4305
rect 17645 4225 17665 4305
rect 17735 4225 17755 4305
rect 17825 4225 17845 4305
rect 17915 4225 17935 4305
rect 18005 4225 18025 4305
rect 18095 4225 18115 4305
rect 18185 4225 18205 4305
rect 18275 4225 18295 4305
rect 18365 4225 18385 4305
rect 18455 4225 18475 4305
rect 18545 4225 18565 4305
rect 18635 4225 18655 4305
rect 18725 4225 18745 4305
rect 18815 4225 18835 4305
rect 18905 4225 18925 4305
rect 18995 4225 19015 4305
rect 19085 4225 19105 4305
rect 19175 4225 19195 4305
rect 19265 4225 19285 4305
rect 19355 4225 19375 4305
rect 19445 4225 19465 4305
rect 19535 4225 19555 4305
rect 19625 4225 19645 4305
rect 19715 4225 19735 4305
rect 19805 4225 19825 4305
rect 19895 4225 19915 4305
rect 19985 4225 20005 4305
rect 20705 4225 20725 4305
rect 9950 4170 9970 4190
rect 10130 4170 10150 4190
rect 10310 4170 10330 4190
rect 10490 4170 10510 4190
rect 10670 4170 10690 4190
rect 10850 4170 10870 4190
rect 11030 4170 11050 4190
rect 11210 4170 11230 4190
rect 11390 4170 11410 4190
rect 11570 4170 11590 4190
rect 11750 4170 11770 4190
rect 11930 4170 11950 4190
rect 12110 4170 12130 4190
rect 12290 4170 12310 4190
rect 12470 4170 12490 4190
rect 12650 4170 12670 4190
rect 12830 4170 12850 4190
rect 13010 4170 13030 4190
rect 13190 4170 13210 4190
rect 13370 4170 13390 4190
rect 13550 4170 13570 4190
rect 13730 4170 13750 4190
rect 13910 4170 13930 4190
rect 14090 4170 14110 4190
rect 14270 4170 14290 4190
rect 14450 4170 14470 4190
rect 14630 4170 14650 4190
rect 14810 4170 14830 4190
rect 15080 4170 15100 4190
rect 15260 4170 15280 4190
rect 15440 4170 15460 4190
rect 15620 4170 15640 4190
rect 15800 4170 15820 4190
rect 15980 4170 16000 4190
rect 16160 4170 16180 4190
rect 16340 4170 16360 4190
rect 16520 4170 16540 4190
rect 16700 4170 16720 4190
rect 16880 4170 16900 4190
rect 17060 4170 17080 4190
rect 17240 4170 17260 4190
rect 17420 4170 17440 4190
rect 17600 4170 17620 4190
rect 17780 4170 17800 4190
rect 17960 4170 17980 4190
rect 18140 4170 18160 4190
rect 18320 4170 18340 4190
rect 18500 4170 18520 4190
rect 18680 4170 18700 4190
rect 18860 4170 18880 4190
rect 19040 4170 19060 4190
rect 19220 4170 19240 4190
rect 19400 4170 19420 4190
rect 19580 4170 19600 4190
rect 19760 4170 19780 4190
rect 19940 4170 19960 4190
rect 10040 4085 10060 4105
rect 10580 4085 10600 4105
rect 10760 4085 10780 4105
rect 11300 4085 11320 4105
rect 11480 4085 11500 4105
rect 12020 4085 12040 4105
rect 12200 4085 12220 4105
rect 12740 4085 12760 4105
rect 12920 4085 12940 4105
rect 13460 4085 13480 4105
rect 13640 4085 13660 4105
rect 13775 4085 13795 4105
rect 13865 4085 13885 4105
rect 13955 4085 13975 4105
rect 14180 4085 14200 4105
rect 15710 4085 15730 4105
rect 15935 4085 15955 4105
rect 16025 4085 16045 4105
rect 16115 4085 16135 4105
rect 16250 4085 16270 4105
rect 16430 4085 16450 4105
rect 16970 4085 16990 4105
rect 17150 4085 17170 4105
rect 17690 4085 17710 4105
rect 17870 4085 17890 4105
rect 18410 4085 18430 4105
rect 18590 4085 18610 4105
rect 19130 4085 19150 4105
rect 19310 4085 19330 4105
rect 19850 4085 19870 4105
rect 13550 4005 13570 4025
rect 14090 4005 14110 4025
rect 15800 4005 15820 4025
rect 16340 4005 16360 4025
rect 20345 4005 20365 4025
rect 13730 3965 13750 3985
rect 13910 3965 13930 3985
rect 15980 3965 16000 3985
rect 16160 3965 16180 3985
rect 20435 3965 20455 3985
rect 10085 3925 10105 3945
rect 10265 3925 10285 3945
rect 10445 3925 10465 3945
rect 10805 3925 10825 3945
rect 10985 3925 11005 3945
rect 11165 3925 11185 3945
rect 11525 3925 11545 3945
rect 11705 3925 11725 3945
rect 11885 3925 11905 3945
rect 12245 3925 12265 3945
rect 12425 3925 12445 3945
rect 12605 3925 12625 3945
rect 12965 3925 12985 3945
rect 13145 3925 13165 3945
rect 13325 3925 13345 3945
rect 14405 3925 14425 3945
rect 14585 3925 14605 3945
rect 14765 3925 14785 3945
rect 15125 3925 15145 3945
rect 15305 3925 15325 3945
rect 15485 3925 15505 3945
rect 16565 3925 16585 3945
rect 16745 3925 16765 3945
rect 16925 3925 16945 3945
rect 17285 3925 17305 3945
rect 17465 3925 17485 3945
rect 17645 3925 17665 3945
rect 18005 3925 18025 3945
rect 18185 3925 18205 3945
rect 18365 3925 18385 3945
rect 18725 3925 18745 3945
rect 18905 3925 18925 3945
rect 19085 3925 19105 3945
rect 19445 3925 19465 3945
rect 19625 3925 19645 3945
rect 19805 3925 19825 3945
rect 10130 3885 10150 3905
rect 10175 3885 10195 3905
rect 10220 3885 10240 3905
rect 10310 3885 10330 3905
rect 10355 3885 10375 3905
rect 10400 3885 10420 3905
rect 10850 3885 10870 3905
rect 10895 3885 10915 3905
rect 10940 3885 10960 3905
rect 11030 3885 11050 3905
rect 11075 3885 11095 3905
rect 11120 3885 11140 3905
rect 11570 3885 11590 3905
rect 11615 3885 11635 3905
rect 11660 3885 11680 3905
rect 11750 3885 11770 3905
rect 11795 3885 11815 3905
rect 11840 3885 11860 3905
rect 12290 3885 12310 3905
rect 12335 3885 12355 3905
rect 12380 3885 12400 3905
rect 12470 3885 12490 3905
rect 12515 3885 12535 3905
rect 12560 3885 12580 3905
rect 13010 3885 13030 3905
rect 13055 3885 13075 3905
rect 13100 3885 13120 3905
rect 13190 3885 13210 3905
rect 13235 3885 13255 3905
rect 13280 3885 13300 3905
rect 16610 3885 16630 3905
rect 16655 3885 16675 3905
rect 16700 3885 16720 3905
rect 16790 3885 16810 3905
rect 16835 3885 16855 3905
rect 16880 3885 16900 3905
rect 17330 3885 17350 3905
rect 17375 3885 17395 3905
rect 17420 3885 17440 3905
rect 17510 3885 17530 3905
rect 17555 3885 17575 3905
rect 17600 3885 17620 3905
rect 18050 3885 18070 3905
rect 18095 3885 18115 3905
rect 18140 3885 18160 3905
rect 18230 3885 18250 3905
rect 18275 3885 18295 3905
rect 18320 3885 18340 3905
rect 18770 3885 18790 3905
rect 18815 3885 18835 3905
rect 18860 3885 18880 3905
rect 18950 3885 18970 3905
rect 18995 3885 19015 3905
rect 19040 3885 19060 3905
rect 19490 3885 19510 3905
rect 19535 3885 19555 3905
rect 19580 3885 19600 3905
rect 19670 3885 19690 3905
rect 19715 3885 19735 3905
rect 19760 3885 19780 3905
rect 13820 3845 13840 3865
rect 14000 3845 14020 3865
rect 14450 3845 14470 3865
rect 14630 3845 14650 3865
rect 15260 3845 15280 3865
rect 15440 3845 15460 3865
rect 15890 3845 15910 3865
rect 16070 3845 16090 3865
rect 10085 3805 10105 3825
rect 10265 3805 10285 3825
rect 10445 3805 10465 3825
rect 10805 3805 10825 3825
rect 10985 3805 11005 3825
rect 11165 3805 11185 3825
rect 11525 3805 11545 3825
rect 11705 3805 11725 3825
rect 11885 3805 11905 3825
rect 12245 3805 12265 3825
rect 12425 3805 12445 3825
rect 12605 3805 12625 3825
rect 12965 3805 12985 3825
rect 13145 3805 13165 3825
rect 13325 3805 13345 3825
rect 13685 3805 13705 3825
rect 13865 3805 13885 3825
rect 14045 3805 14065 3825
rect 15845 3805 15865 3825
rect 16025 3805 16045 3825
rect 16205 3805 16225 3825
rect 16565 3805 16585 3825
rect 16745 3805 16765 3825
rect 16925 3805 16945 3825
rect 17285 3805 17305 3825
rect 17465 3805 17485 3825
rect 17645 3805 17665 3825
rect 18005 3805 18025 3825
rect 18185 3805 18205 3825
rect 18365 3805 18385 3825
rect 18725 3805 18745 3825
rect 18905 3805 18925 3825
rect 19085 3805 19105 3825
rect 19445 3805 19465 3825
rect 19625 3805 19645 3825
rect 19805 3805 19825 3825
rect 9950 3765 9970 3785
rect 10490 3765 10510 3785
rect 10670 3765 10690 3785
rect 11210 3765 11230 3785
rect 11390 3765 11410 3785
rect 11930 3765 11950 3785
rect 12110 3765 12130 3785
rect 12650 3765 12670 3785
rect 12830 3765 12850 3785
rect 13370 3765 13390 3785
rect 14270 3765 14290 3785
rect 14495 3765 14515 3785
rect 14585 3765 14605 3785
rect 14675 3765 14695 3785
rect 14810 3765 14830 3785
rect 15080 3765 15100 3785
rect 15215 3765 15235 3785
rect 15305 3765 15325 3785
rect 15395 3765 15415 3785
rect 15620 3765 15640 3785
rect 16520 3765 16540 3785
rect 17060 3765 17080 3785
rect 17240 3765 17260 3785
rect 17780 3765 17800 3785
rect 17960 3765 17980 3785
rect 18500 3765 18520 3785
rect 18680 3765 18700 3785
rect 19220 3765 19240 3785
rect 19400 3765 19420 3785
rect 19940 3765 19960 3785
rect 14540 3725 14560 3745
rect 14720 3725 14740 3745
rect 15170 3725 15190 3745
rect 15350 3725 15370 3745
rect 20615 3725 20635 3745
rect 14360 3685 14380 3705
rect 14900 3685 14920 3705
rect 14990 3685 15010 3705
rect 15530 3685 15550 3705
rect 20525 3685 20545 3705
rect 10040 3600 10060 3620
rect 10220 3600 10240 3620
rect 10400 3600 10420 3620
rect 10580 3600 10600 3620
rect 10760 3600 10780 3620
rect 10940 3600 10960 3620
rect 11120 3600 11140 3620
rect 11300 3600 11320 3620
rect 11480 3600 11500 3620
rect 11660 3600 11680 3620
rect 11840 3600 11860 3620
rect 12020 3600 12040 3620
rect 12200 3600 12220 3620
rect 12380 3600 12400 3620
rect 12560 3600 12580 3620
rect 12740 3600 12760 3620
rect 12920 3600 12940 3620
rect 13100 3600 13120 3620
rect 13280 3600 13300 3620
rect 13460 3600 13480 3620
rect 13640 3600 13660 3620
rect 13820 3600 13840 3620
rect 14000 3600 14020 3620
rect 14180 3600 14200 3620
rect 14360 3600 14380 3620
rect 14540 3600 14560 3620
rect 14720 3600 14740 3620
rect 14900 3600 14920 3620
rect 14990 3600 15010 3620
rect 15170 3600 15190 3620
rect 15350 3600 15370 3620
rect 15530 3600 15550 3620
rect 15710 3600 15730 3620
rect 15890 3600 15910 3620
rect 16070 3600 16090 3620
rect 16250 3600 16270 3620
rect 16430 3600 16450 3620
rect 16610 3600 16630 3620
rect 16790 3600 16810 3620
rect 16970 3600 16990 3620
rect 17150 3600 17170 3620
rect 17330 3600 17350 3620
rect 17510 3600 17530 3620
rect 17690 3600 17710 3620
rect 17870 3600 17890 3620
rect 18050 3600 18070 3620
rect 18230 3600 18250 3620
rect 18410 3600 18430 3620
rect 18590 3600 18610 3620
rect 18770 3600 18790 3620
rect 18950 3600 18970 3620
rect 19130 3600 19150 3620
rect 19310 3600 19330 3620
rect 19490 3600 19510 3620
rect 19670 3600 19690 3620
rect 19850 3600 19870 3620
rect 9185 3485 9205 3565
rect 9905 3485 9925 3565
rect 9995 3485 10015 3565
rect 10085 3485 10105 3565
rect 10175 3485 10195 3565
rect 10265 3485 10285 3565
rect 10355 3485 10375 3565
rect 10445 3485 10465 3565
rect 10535 3485 10555 3565
rect 10625 3485 10645 3565
rect 10715 3485 10735 3565
rect 10805 3485 10825 3565
rect 10895 3485 10915 3565
rect 10985 3485 11005 3565
rect 11075 3485 11095 3565
rect 11165 3485 11185 3565
rect 11255 3485 11275 3565
rect 11345 3485 11365 3565
rect 11435 3485 11455 3565
rect 11525 3485 11545 3565
rect 11615 3485 11635 3565
rect 11705 3485 11725 3565
rect 11795 3485 11815 3565
rect 11885 3485 11905 3565
rect 11975 3485 11995 3565
rect 12065 3485 12085 3565
rect 12155 3485 12175 3565
rect 12245 3485 12265 3565
rect 12335 3485 12355 3565
rect 12425 3485 12445 3565
rect 12515 3485 12535 3565
rect 12605 3485 12625 3565
rect 12695 3485 12715 3565
rect 12785 3485 12805 3565
rect 12875 3485 12895 3565
rect 12965 3485 12985 3565
rect 13055 3485 13075 3565
rect 13145 3485 13165 3565
rect 13235 3485 13255 3565
rect 13325 3485 13345 3565
rect 13415 3485 13435 3565
rect 13505 3485 13525 3565
rect 13595 3485 13615 3565
rect 13685 3485 13705 3565
rect 13775 3485 13795 3565
rect 13865 3485 13885 3565
rect 13955 3485 13975 3565
rect 14045 3485 14065 3565
rect 14135 3485 14155 3565
rect 14225 3485 14245 3565
rect 14315 3485 14335 3565
rect 14405 3485 14425 3565
rect 14495 3485 14515 3565
rect 14585 3485 14605 3565
rect 14675 3485 14695 3565
rect 14765 3485 14785 3565
rect 14855 3485 14875 3565
rect 14945 3485 14965 3565
rect 15035 3485 15055 3565
rect 15125 3485 15145 3565
rect 15215 3485 15235 3565
rect 15305 3485 15325 3565
rect 15395 3485 15415 3565
rect 15485 3485 15505 3565
rect 15575 3485 15595 3565
rect 15665 3485 15685 3565
rect 15755 3485 15775 3565
rect 15845 3485 15865 3565
rect 15935 3485 15955 3565
rect 16025 3485 16045 3565
rect 16115 3485 16135 3565
rect 16205 3485 16225 3565
rect 16295 3485 16315 3565
rect 16385 3485 16405 3565
rect 16475 3485 16495 3565
rect 16565 3485 16585 3565
rect 16655 3485 16675 3565
rect 16745 3485 16765 3565
rect 16835 3485 16855 3565
rect 16925 3485 16945 3565
rect 17015 3485 17035 3565
rect 17105 3485 17125 3565
rect 17195 3485 17215 3565
rect 17285 3485 17305 3565
rect 17375 3485 17395 3565
rect 17465 3485 17485 3565
rect 17555 3485 17575 3565
rect 17645 3485 17665 3565
rect 17735 3485 17755 3565
rect 17825 3485 17845 3565
rect 17915 3485 17935 3565
rect 18005 3485 18025 3565
rect 18095 3485 18115 3565
rect 18185 3485 18205 3565
rect 18275 3485 18295 3565
rect 18365 3485 18385 3565
rect 18455 3485 18475 3565
rect 18545 3485 18565 3565
rect 18635 3485 18655 3565
rect 18725 3485 18745 3565
rect 18815 3485 18835 3565
rect 18905 3485 18925 3565
rect 18995 3485 19015 3565
rect 19085 3485 19105 3565
rect 19175 3485 19195 3565
rect 19265 3485 19285 3565
rect 19355 3485 19375 3565
rect 19445 3485 19465 3565
rect 19535 3485 19555 3565
rect 19625 3485 19645 3565
rect 19715 3485 19735 3565
rect 19805 3485 19825 3565
rect 19895 3485 19915 3565
rect 19985 3485 20005 3565
rect 20705 3485 20725 3565
rect 9050 3425 9070 3445
rect 9185 3425 9205 3445
rect 9905 3425 9925 3445
rect 10085 3425 10105 3445
rect 10265 3425 10285 3445
rect 10445 3425 10465 3445
rect 10625 3425 10645 3445
rect 10805 3425 10825 3445
rect 10985 3425 11005 3445
rect 11165 3425 11185 3445
rect 11345 3425 11365 3445
rect 11525 3425 11545 3445
rect 11705 3425 11725 3445
rect 11885 3425 11905 3445
rect 12065 3425 12085 3445
rect 12245 3425 12265 3445
rect 12425 3425 12445 3445
rect 12605 3425 12625 3445
rect 12785 3425 12805 3445
rect 12965 3425 12985 3445
rect 13145 3425 13165 3445
rect 13325 3425 13345 3445
rect 13505 3425 13525 3445
rect 13685 3425 13705 3445
rect 13865 3425 13885 3445
rect 14045 3425 14065 3445
rect 14225 3425 14245 3445
rect 14405 3425 14425 3445
rect 14585 3425 14605 3445
rect 14765 3425 14785 3445
rect 14945 3425 14965 3445
rect 15125 3425 15145 3445
rect 15305 3425 15325 3445
rect 15485 3425 15505 3445
rect 15665 3425 15685 3445
rect 15845 3425 15865 3445
rect 16025 3425 16045 3445
rect 16205 3425 16225 3445
rect 16385 3425 16405 3445
rect 16565 3425 16585 3445
rect 16745 3425 16765 3445
rect 16925 3425 16945 3445
rect 17105 3425 17125 3445
rect 17285 3425 17305 3445
rect 17465 3425 17485 3445
rect 17645 3425 17665 3445
rect 17825 3425 17845 3445
rect 18005 3425 18025 3445
rect 18185 3425 18205 3445
rect 18365 3425 18385 3445
rect 18545 3425 18565 3445
rect 18725 3425 18745 3445
rect 18905 3425 18925 3445
rect 19085 3425 19105 3445
rect 19265 3425 19285 3445
rect 19445 3425 19465 3445
rect 19625 3425 19645 3445
rect 19805 3425 19825 3445
rect 19985 3425 20005 3445
rect 20705 3425 20725 3445
rect 20840 3425 20860 3445
<< metal1 >>
rect 9040 3450 9080 4375
rect 9175 4370 9215 4375
rect 9175 4340 9180 4370
rect 9210 4340 9215 4370
rect 9175 4335 9215 4340
rect 9185 4315 9205 4335
rect 9275 4315 9295 4375
rect 9365 4315 9385 4375
rect 9455 4315 9475 4375
rect 9545 4315 9565 4375
rect 9635 4315 9655 4375
rect 9725 4315 9745 4375
rect 9815 4315 9835 4375
rect 9895 4370 9935 4375
rect 9895 4340 9900 4370
rect 9930 4340 9935 4370
rect 9895 4335 9935 4340
rect 10075 4370 10115 4375
rect 10075 4340 10080 4370
rect 10110 4340 10115 4370
rect 10075 4335 10115 4340
rect 10255 4370 10295 4375
rect 10255 4340 10260 4370
rect 10290 4340 10295 4370
rect 10255 4335 10295 4340
rect 10435 4370 10475 4375
rect 10435 4340 10440 4370
rect 10470 4340 10475 4370
rect 10435 4335 10475 4340
rect 10615 4370 10655 4375
rect 10615 4340 10620 4370
rect 10650 4340 10655 4370
rect 10615 4335 10655 4340
rect 10795 4370 10835 4375
rect 10795 4340 10800 4370
rect 10830 4340 10835 4370
rect 10795 4335 10835 4340
rect 10975 4370 11015 4375
rect 10975 4340 10980 4370
rect 11010 4340 11015 4370
rect 10975 4335 11015 4340
rect 11155 4370 11195 4375
rect 11155 4340 11160 4370
rect 11190 4340 11195 4370
rect 11155 4335 11195 4340
rect 11335 4370 11375 4375
rect 11335 4340 11340 4370
rect 11370 4340 11375 4370
rect 11335 4335 11375 4340
rect 11515 4370 11555 4375
rect 11515 4340 11520 4370
rect 11550 4340 11555 4370
rect 11515 4335 11555 4340
rect 11695 4370 11735 4375
rect 11695 4340 11700 4370
rect 11730 4340 11735 4370
rect 11695 4335 11735 4340
rect 11875 4370 11915 4375
rect 11875 4340 11880 4370
rect 11910 4340 11915 4370
rect 11875 4335 11915 4340
rect 12055 4370 12095 4375
rect 12055 4340 12060 4370
rect 12090 4340 12095 4370
rect 12055 4335 12095 4340
rect 12235 4370 12275 4375
rect 12235 4340 12240 4370
rect 12270 4340 12275 4370
rect 12235 4335 12275 4340
rect 12415 4370 12455 4375
rect 12415 4340 12420 4370
rect 12450 4340 12455 4370
rect 12415 4335 12455 4340
rect 12595 4370 12635 4375
rect 12595 4340 12600 4370
rect 12630 4340 12635 4370
rect 12595 4335 12635 4340
rect 12775 4370 12815 4375
rect 12775 4340 12780 4370
rect 12810 4340 12815 4370
rect 12775 4335 12815 4340
rect 12955 4370 12995 4375
rect 12955 4340 12960 4370
rect 12990 4340 12995 4370
rect 12955 4335 12995 4340
rect 13135 4370 13175 4375
rect 13135 4340 13140 4370
rect 13170 4340 13175 4370
rect 13135 4335 13175 4340
rect 13315 4370 13355 4375
rect 13315 4340 13320 4370
rect 13350 4340 13355 4370
rect 13315 4335 13355 4340
rect 13495 4370 13535 4375
rect 13495 4340 13500 4370
rect 13530 4340 13535 4370
rect 13495 4335 13535 4340
rect 13675 4370 13715 4375
rect 13675 4340 13680 4370
rect 13710 4340 13715 4370
rect 13675 4335 13715 4340
rect 13855 4370 13895 4375
rect 13855 4340 13860 4370
rect 13890 4340 13895 4370
rect 13855 4335 13895 4340
rect 14035 4370 14075 4375
rect 14035 4340 14040 4370
rect 14070 4340 14075 4370
rect 14035 4335 14075 4340
rect 14215 4370 14255 4375
rect 14215 4340 14220 4370
rect 14250 4340 14255 4370
rect 14215 4335 14255 4340
rect 14395 4370 14435 4375
rect 14395 4340 14400 4370
rect 14430 4340 14435 4370
rect 14395 4335 14435 4340
rect 14575 4370 14615 4375
rect 14575 4340 14580 4370
rect 14610 4340 14615 4370
rect 14575 4335 14615 4340
rect 14755 4370 14795 4375
rect 14755 4340 14760 4370
rect 14790 4340 14795 4370
rect 14755 4335 14795 4340
rect 14935 4370 14975 4375
rect 14935 4340 14940 4370
rect 14970 4340 14975 4370
rect 14935 4335 14975 4340
rect 15115 4370 15155 4375
rect 15115 4340 15120 4370
rect 15150 4340 15155 4370
rect 15115 4335 15155 4340
rect 15295 4370 15335 4375
rect 15295 4340 15300 4370
rect 15330 4340 15335 4370
rect 15295 4335 15335 4340
rect 15475 4370 15515 4375
rect 15475 4340 15480 4370
rect 15510 4340 15515 4370
rect 15475 4335 15515 4340
rect 15655 4370 15695 4375
rect 15655 4340 15660 4370
rect 15690 4340 15695 4370
rect 15655 4335 15695 4340
rect 15835 4370 15875 4375
rect 15835 4340 15840 4370
rect 15870 4340 15875 4370
rect 15835 4335 15875 4340
rect 16015 4370 16055 4375
rect 16015 4340 16020 4370
rect 16050 4340 16055 4370
rect 16015 4335 16055 4340
rect 16195 4370 16235 4375
rect 16195 4340 16200 4370
rect 16230 4340 16235 4370
rect 16195 4335 16235 4340
rect 16375 4370 16415 4375
rect 16375 4340 16380 4370
rect 16410 4340 16415 4370
rect 16375 4335 16415 4340
rect 16555 4370 16595 4375
rect 16555 4340 16560 4370
rect 16590 4340 16595 4370
rect 16555 4335 16595 4340
rect 16735 4370 16775 4375
rect 16735 4340 16740 4370
rect 16770 4340 16775 4370
rect 16735 4335 16775 4340
rect 16915 4370 16955 4375
rect 16915 4340 16920 4370
rect 16950 4340 16955 4370
rect 16915 4335 16955 4340
rect 17095 4370 17135 4375
rect 17095 4340 17100 4370
rect 17130 4340 17135 4370
rect 17095 4335 17135 4340
rect 17275 4370 17315 4375
rect 17275 4340 17280 4370
rect 17310 4340 17315 4370
rect 17275 4335 17315 4340
rect 17455 4370 17495 4375
rect 17455 4340 17460 4370
rect 17490 4340 17495 4370
rect 17455 4335 17495 4340
rect 17635 4370 17675 4375
rect 17635 4340 17640 4370
rect 17670 4340 17675 4370
rect 17635 4335 17675 4340
rect 17815 4370 17855 4375
rect 17815 4340 17820 4370
rect 17850 4340 17855 4370
rect 17815 4335 17855 4340
rect 17995 4370 18035 4375
rect 17995 4340 18000 4370
rect 18030 4340 18035 4370
rect 17995 4335 18035 4340
rect 18175 4370 18215 4375
rect 18175 4340 18180 4370
rect 18210 4340 18215 4370
rect 18175 4335 18215 4340
rect 18355 4370 18395 4375
rect 18355 4340 18360 4370
rect 18390 4340 18395 4370
rect 18355 4335 18395 4340
rect 18535 4370 18575 4375
rect 18535 4340 18540 4370
rect 18570 4340 18575 4370
rect 18535 4335 18575 4340
rect 18715 4370 18755 4375
rect 18715 4340 18720 4370
rect 18750 4340 18755 4370
rect 18715 4335 18755 4340
rect 18895 4370 18935 4375
rect 18895 4340 18900 4370
rect 18930 4340 18935 4370
rect 18895 4335 18935 4340
rect 19075 4370 19115 4375
rect 19075 4340 19080 4370
rect 19110 4340 19115 4370
rect 19075 4335 19115 4340
rect 19255 4370 19295 4375
rect 19255 4340 19260 4370
rect 19290 4340 19295 4370
rect 19255 4335 19295 4340
rect 19435 4370 19475 4375
rect 19435 4340 19440 4370
rect 19470 4340 19475 4370
rect 19435 4335 19475 4340
rect 19615 4370 19655 4375
rect 19615 4340 19620 4370
rect 19650 4340 19655 4370
rect 19615 4335 19655 4340
rect 19795 4370 19835 4375
rect 19795 4340 19800 4370
rect 19830 4340 19835 4370
rect 19795 4335 19835 4340
rect 19975 4370 20015 4375
rect 19975 4340 19980 4370
rect 20010 4340 20015 4370
rect 19975 4335 20015 4340
rect 9905 4315 9925 4335
rect 10625 4315 10645 4335
rect 11345 4315 11365 4335
rect 12065 4315 12085 4335
rect 12785 4315 12805 4335
rect 13505 4315 13525 4335
rect 14225 4315 14245 4335
rect 14945 4315 14965 4335
rect 15665 4315 15685 4335
rect 16385 4315 16405 4335
rect 17105 4315 17125 4335
rect 17825 4315 17845 4335
rect 18545 4315 18565 4335
rect 19265 4315 19285 4335
rect 19985 4315 20005 4335
rect 20075 4315 20095 4375
rect 20165 4315 20185 4375
rect 20255 4315 20275 4375
rect 20345 4315 20365 4375
rect 20435 4315 20455 4375
rect 20525 4315 20545 4375
rect 20615 4315 20635 4375
rect 20695 4370 20735 4375
rect 20695 4340 20700 4370
rect 20730 4340 20735 4370
rect 20695 4335 20735 4340
rect 20705 4315 20725 4335
rect 9180 4305 9210 4315
rect 9180 4225 9185 4305
rect 9205 4225 9210 4305
rect 9180 4215 9210 4225
rect 9270 4215 9300 4315
rect 9360 4215 9390 4315
rect 9450 4215 9480 4315
rect 9540 4215 9570 4315
rect 9630 4215 9660 4315
rect 9720 4215 9750 4315
rect 9810 4215 9840 4315
rect 9900 4305 9930 4315
rect 9900 4225 9905 4305
rect 9925 4225 9930 4305
rect 9900 4215 9930 4225
rect 9990 4305 10020 4315
rect 9990 4225 9995 4305
rect 10015 4225 10020 4305
rect 9990 4215 10020 4225
rect 10080 4305 10110 4315
rect 10080 4225 10085 4305
rect 10105 4225 10110 4305
rect 10080 4215 10110 4225
rect 10170 4305 10200 4315
rect 10170 4225 10175 4305
rect 10195 4225 10200 4305
rect 10170 4215 10200 4225
rect 10260 4305 10290 4315
rect 10260 4225 10265 4305
rect 10285 4225 10290 4305
rect 10260 4215 10290 4225
rect 10350 4305 10380 4315
rect 10350 4225 10355 4305
rect 10375 4225 10380 4305
rect 10350 4215 10380 4225
rect 10440 4305 10470 4315
rect 10440 4225 10445 4305
rect 10465 4225 10470 4305
rect 10440 4215 10470 4225
rect 10530 4305 10560 4315
rect 10530 4225 10535 4305
rect 10555 4225 10560 4305
rect 10530 4215 10560 4225
rect 10620 4305 10650 4315
rect 10620 4225 10625 4305
rect 10645 4225 10650 4305
rect 10620 4215 10650 4225
rect 10710 4305 10740 4315
rect 10710 4225 10715 4305
rect 10735 4225 10740 4305
rect 10710 4215 10740 4225
rect 10800 4305 10830 4315
rect 10800 4225 10805 4305
rect 10825 4225 10830 4305
rect 10800 4215 10830 4225
rect 10890 4305 10920 4315
rect 10890 4225 10895 4305
rect 10915 4225 10920 4305
rect 10890 4215 10920 4225
rect 10980 4305 11010 4315
rect 10980 4225 10985 4305
rect 11005 4225 11010 4305
rect 10980 4215 11010 4225
rect 11070 4305 11100 4315
rect 11070 4225 11075 4305
rect 11095 4225 11100 4305
rect 11070 4215 11100 4225
rect 11160 4305 11190 4315
rect 11160 4225 11165 4305
rect 11185 4225 11190 4305
rect 11160 4215 11190 4225
rect 11250 4305 11280 4315
rect 11250 4225 11255 4305
rect 11275 4225 11280 4305
rect 11250 4215 11280 4225
rect 11340 4305 11370 4315
rect 11340 4225 11345 4305
rect 11365 4225 11370 4305
rect 11340 4215 11370 4225
rect 11430 4305 11460 4315
rect 11430 4225 11435 4305
rect 11455 4225 11460 4305
rect 11430 4215 11460 4225
rect 11520 4305 11550 4315
rect 11520 4225 11525 4305
rect 11545 4225 11550 4305
rect 11520 4215 11550 4225
rect 11610 4305 11640 4315
rect 11610 4225 11615 4305
rect 11635 4225 11640 4305
rect 11610 4215 11640 4225
rect 11700 4305 11730 4315
rect 11700 4225 11705 4305
rect 11725 4225 11730 4305
rect 11700 4215 11730 4225
rect 11790 4305 11820 4315
rect 11790 4225 11795 4305
rect 11815 4225 11820 4305
rect 11790 4215 11820 4225
rect 11880 4305 11910 4315
rect 11880 4225 11885 4305
rect 11905 4225 11910 4305
rect 11880 4215 11910 4225
rect 11970 4305 12000 4315
rect 11970 4225 11975 4305
rect 11995 4225 12000 4305
rect 11970 4215 12000 4225
rect 12060 4305 12090 4315
rect 12060 4225 12065 4305
rect 12085 4225 12090 4305
rect 12060 4215 12090 4225
rect 12150 4305 12180 4315
rect 12150 4225 12155 4305
rect 12175 4225 12180 4305
rect 12150 4215 12180 4225
rect 12240 4305 12270 4315
rect 12240 4225 12245 4305
rect 12265 4225 12270 4305
rect 12240 4215 12270 4225
rect 12330 4305 12360 4315
rect 12330 4225 12335 4305
rect 12355 4225 12360 4305
rect 12330 4215 12360 4225
rect 12420 4305 12450 4315
rect 12420 4225 12425 4305
rect 12445 4225 12450 4305
rect 12420 4215 12450 4225
rect 12510 4305 12540 4315
rect 12510 4225 12515 4305
rect 12535 4225 12540 4305
rect 12510 4215 12540 4225
rect 12600 4305 12630 4315
rect 12600 4225 12605 4305
rect 12625 4225 12630 4305
rect 12600 4215 12630 4225
rect 12690 4305 12720 4315
rect 12690 4225 12695 4305
rect 12715 4225 12720 4305
rect 12690 4215 12720 4225
rect 12780 4305 12810 4315
rect 12780 4225 12785 4305
rect 12805 4225 12810 4305
rect 12780 4215 12810 4225
rect 12870 4305 12900 4315
rect 12870 4225 12875 4305
rect 12895 4225 12900 4305
rect 12870 4215 12900 4225
rect 12960 4305 12990 4315
rect 12960 4225 12965 4305
rect 12985 4225 12990 4305
rect 12960 4215 12990 4225
rect 13050 4305 13080 4315
rect 13050 4225 13055 4305
rect 13075 4225 13080 4305
rect 13050 4215 13080 4225
rect 13140 4305 13170 4315
rect 13140 4225 13145 4305
rect 13165 4225 13170 4305
rect 13140 4215 13170 4225
rect 13230 4305 13260 4315
rect 13230 4225 13235 4305
rect 13255 4225 13260 4305
rect 13230 4215 13260 4225
rect 13320 4305 13350 4315
rect 13320 4225 13325 4305
rect 13345 4225 13350 4305
rect 13320 4215 13350 4225
rect 13410 4305 13440 4315
rect 13410 4225 13415 4305
rect 13435 4225 13440 4305
rect 13410 4215 13440 4225
rect 13500 4305 13530 4315
rect 13500 4225 13505 4305
rect 13525 4225 13530 4305
rect 13500 4215 13530 4225
rect 13590 4305 13620 4315
rect 13590 4225 13595 4305
rect 13615 4225 13620 4305
rect 13590 4215 13620 4225
rect 13680 4305 13710 4315
rect 13680 4225 13685 4305
rect 13705 4225 13710 4305
rect 13680 4215 13710 4225
rect 13770 4305 13800 4315
rect 13770 4225 13775 4305
rect 13795 4225 13800 4305
rect 13770 4215 13800 4225
rect 13860 4305 13890 4315
rect 13860 4225 13865 4305
rect 13885 4225 13890 4305
rect 13860 4215 13890 4225
rect 13950 4305 13980 4315
rect 13950 4225 13955 4305
rect 13975 4225 13980 4305
rect 13950 4215 13980 4225
rect 14040 4305 14070 4315
rect 14040 4225 14045 4305
rect 14065 4225 14070 4305
rect 14040 4215 14070 4225
rect 14130 4305 14160 4315
rect 14130 4225 14135 4305
rect 14155 4225 14160 4305
rect 14130 4215 14160 4225
rect 14220 4305 14250 4315
rect 14220 4225 14225 4305
rect 14245 4225 14250 4305
rect 14220 4215 14250 4225
rect 14310 4305 14340 4315
rect 14310 4225 14315 4305
rect 14335 4225 14340 4305
rect 14310 4215 14340 4225
rect 14400 4305 14430 4315
rect 14400 4225 14405 4305
rect 14425 4225 14430 4305
rect 14400 4215 14430 4225
rect 14490 4305 14520 4315
rect 14490 4225 14495 4305
rect 14515 4225 14520 4305
rect 14490 4215 14520 4225
rect 14580 4305 14610 4315
rect 14580 4225 14585 4305
rect 14605 4225 14610 4305
rect 14580 4215 14610 4225
rect 14670 4305 14700 4315
rect 14670 4225 14675 4305
rect 14695 4225 14700 4305
rect 14670 4215 14700 4225
rect 14760 4305 14790 4315
rect 14760 4225 14765 4305
rect 14785 4225 14790 4305
rect 14760 4215 14790 4225
rect 14850 4305 14880 4315
rect 14850 4225 14855 4305
rect 14875 4225 14880 4305
rect 14850 4215 14880 4225
rect 14940 4305 14970 4315
rect 14940 4225 14945 4305
rect 14965 4225 14970 4305
rect 14940 4215 14970 4225
rect 15030 4305 15060 4315
rect 15030 4225 15035 4305
rect 15055 4225 15060 4305
rect 15030 4215 15060 4225
rect 15120 4305 15150 4315
rect 15120 4225 15125 4305
rect 15145 4225 15150 4305
rect 15120 4215 15150 4225
rect 15210 4305 15240 4315
rect 15210 4225 15215 4305
rect 15235 4225 15240 4305
rect 15210 4215 15240 4225
rect 15300 4305 15330 4315
rect 15300 4225 15305 4305
rect 15325 4225 15330 4305
rect 15300 4215 15330 4225
rect 15390 4305 15420 4315
rect 15390 4225 15395 4305
rect 15415 4225 15420 4305
rect 15390 4215 15420 4225
rect 15480 4305 15510 4315
rect 15480 4225 15485 4305
rect 15505 4225 15510 4305
rect 15480 4215 15510 4225
rect 15570 4305 15600 4315
rect 15570 4225 15575 4305
rect 15595 4225 15600 4305
rect 15570 4215 15600 4225
rect 15660 4305 15690 4315
rect 15660 4225 15665 4305
rect 15685 4225 15690 4305
rect 15660 4215 15690 4225
rect 15750 4305 15780 4315
rect 15750 4225 15755 4305
rect 15775 4225 15780 4305
rect 15750 4215 15780 4225
rect 15840 4305 15870 4315
rect 15840 4225 15845 4305
rect 15865 4225 15870 4305
rect 15840 4215 15870 4225
rect 15930 4305 15960 4315
rect 15930 4225 15935 4305
rect 15955 4225 15960 4305
rect 15930 4215 15960 4225
rect 16020 4305 16050 4315
rect 16020 4225 16025 4305
rect 16045 4225 16050 4305
rect 16020 4215 16050 4225
rect 16110 4305 16140 4315
rect 16110 4225 16115 4305
rect 16135 4225 16140 4305
rect 16110 4215 16140 4225
rect 16200 4305 16230 4315
rect 16200 4225 16205 4305
rect 16225 4225 16230 4305
rect 16200 4215 16230 4225
rect 16290 4305 16320 4315
rect 16290 4225 16295 4305
rect 16315 4225 16320 4305
rect 16290 4215 16320 4225
rect 16380 4305 16410 4315
rect 16380 4225 16385 4305
rect 16405 4225 16410 4305
rect 16380 4215 16410 4225
rect 16470 4305 16500 4315
rect 16470 4225 16475 4305
rect 16495 4225 16500 4305
rect 16470 4215 16500 4225
rect 16560 4305 16590 4315
rect 16560 4225 16565 4305
rect 16585 4225 16590 4305
rect 16560 4215 16590 4225
rect 16650 4305 16680 4315
rect 16650 4225 16655 4305
rect 16675 4225 16680 4305
rect 16650 4215 16680 4225
rect 16740 4305 16770 4315
rect 16740 4225 16745 4305
rect 16765 4225 16770 4305
rect 16740 4215 16770 4225
rect 16830 4305 16860 4315
rect 16830 4225 16835 4305
rect 16855 4225 16860 4305
rect 16830 4215 16860 4225
rect 16920 4305 16950 4315
rect 16920 4225 16925 4305
rect 16945 4225 16950 4305
rect 16920 4215 16950 4225
rect 17010 4305 17040 4315
rect 17010 4225 17015 4305
rect 17035 4225 17040 4305
rect 17010 4215 17040 4225
rect 17100 4305 17130 4315
rect 17100 4225 17105 4305
rect 17125 4225 17130 4305
rect 17100 4215 17130 4225
rect 17190 4305 17220 4315
rect 17190 4225 17195 4305
rect 17215 4225 17220 4305
rect 17190 4215 17220 4225
rect 17280 4305 17310 4315
rect 17280 4225 17285 4305
rect 17305 4225 17310 4305
rect 17280 4215 17310 4225
rect 17370 4305 17400 4315
rect 17370 4225 17375 4305
rect 17395 4225 17400 4305
rect 17370 4215 17400 4225
rect 17460 4305 17490 4315
rect 17460 4225 17465 4305
rect 17485 4225 17490 4305
rect 17460 4215 17490 4225
rect 17550 4305 17580 4315
rect 17550 4225 17555 4305
rect 17575 4225 17580 4305
rect 17550 4215 17580 4225
rect 17640 4305 17670 4315
rect 17640 4225 17645 4305
rect 17665 4225 17670 4305
rect 17640 4215 17670 4225
rect 17730 4305 17760 4315
rect 17730 4225 17735 4305
rect 17755 4225 17760 4305
rect 17730 4215 17760 4225
rect 17820 4305 17850 4315
rect 17820 4225 17825 4305
rect 17845 4225 17850 4305
rect 17820 4215 17850 4225
rect 17910 4305 17940 4315
rect 17910 4225 17915 4305
rect 17935 4225 17940 4305
rect 17910 4215 17940 4225
rect 18000 4305 18030 4315
rect 18000 4225 18005 4305
rect 18025 4225 18030 4305
rect 18000 4215 18030 4225
rect 18090 4305 18120 4315
rect 18090 4225 18095 4305
rect 18115 4225 18120 4305
rect 18090 4215 18120 4225
rect 18180 4305 18210 4315
rect 18180 4225 18185 4305
rect 18205 4225 18210 4305
rect 18180 4215 18210 4225
rect 18270 4305 18300 4315
rect 18270 4225 18275 4305
rect 18295 4225 18300 4305
rect 18270 4215 18300 4225
rect 18360 4305 18390 4315
rect 18360 4225 18365 4305
rect 18385 4225 18390 4305
rect 18360 4215 18390 4225
rect 18450 4305 18480 4315
rect 18450 4225 18455 4305
rect 18475 4225 18480 4305
rect 18450 4215 18480 4225
rect 18540 4305 18570 4315
rect 18540 4225 18545 4305
rect 18565 4225 18570 4305
rect 18540 4215 18570 4225
rect 18630 4305 18660 4315
rect 18630 4225 18635 4305
rect 18655 4225 18660 4305
rect 18630 4215 18660 4225
rect 18720 4305 18750 4315
rect 18720 4225 18725 4305
rect 18745 4225 18750 4305
rect 18720 4215 18750 4225
rect 18810 4305 18840 4315
rect 18810 4225 18815 4305
rect 18835 4225 18840 4305
rect 18810 4215 18840 4225
rect 18900 4305 18930 4315
rect 18900 4225 18905 4305
rect 18925 4225 18930 4305
rect 18900 4215 18930 4225
rect 18990 4305 19020 4315
rect 18990 4225 18995 4305
rect 19015 4225 19020 4305
rect 18990 4215 19020 4225
rect 19080 4305 19110 4315
rect 19080 4225 19085 4305
rect 19105 4225 19110 4305
rect 19080 4215 19110 4225
rect 19170 4305 19200 4315
rect 19170 4225 19175 4305
rect 19195 4225 19200 4305
rect 19170 4215 19200 4225
rect 19260 4305 19290 4315
rect 19260 4225 19265 4305
rect 19285 4225 19290 4305
rect 19260 4215 19290 4225
rect 19350 4305 19380 4315
rect 19350 4225 19355 4305
rect 19375 4225 19380 4305
rect 19350 4215 19380 4225
rect 19440 4305 19470 4315
rect 19440 4225 19445 4305
rect 19465 4225 19470 4305
rect 19440 4215 19470 4225
rect 19530 4305 19560 4315
rect 19530 4225 19535 4305
rect 19555 4225 19560 4305
rect 19530 4215 19560 4225
rect 19620 4305 19650 4315
rect 19620 4225 19625 4305
rect 19645 4225 19650 4305
rect 19620 4215 19650 4225
rect 19710 4305 19740 4315
rect 19710 4225 19715 4305
rect 19735 4225 19740 4305
rect 19710 4215 19740 4225
rect 19800 4305 19830 4315
rect 19800 4225 19805 4305
rect 19825 4225 19830 4305
rect 19800 4215 19830 4225
rect 19890 4305 19920 4315
rect 19890 4225 19895 4305
rect 19915 4225 19920 4305
rect 19890 4215 19920 4225
rect 19980 4305 20010 4315
rect 19980 4225 19985 4305
rect 20005 4225 20010 4305
rect 19980 4215 20010 4225
rect 20070 4215 20100 4315
rect 20160 4215 20190 4315
rect 20250 4215 20280 4315
rect 20340 4215 20370 4315
rect 20430 4215 20460 4315
rect 20520 4215 20550 4315
rect 20610 4215 20640 4315
rect 20700 4305 20730 4315
rect 20700 4225 20705 4305
rect 20725 4225 20730 4305
rect 20700 4215 20730 4225
rect 9275 3575 9295 4215
rect 9365 3575 9385 4215
rect 9455 3575 9475 4215
rect 9545 3575 9565 4215
rect 9635 3575 9655 4215
rect 9725 3575 9745 4215
rect 9815 3575 9835 4215
rect 9950 4195 9970 4200
rect 9945 4190 9975 4195
rect 9945 4170 9950 4190
rect 9970 4170 9975 4190
rect 9945 4165 9975 4170
rect 9950 3790 9970 4165
rect 10040 4110 10060 4115
rect 10035 4105 10065 4110
rect 10035 4085 10040 4105
rect 10060 4085 10065 4105
rect 10035 4080 10065 4085
rect 9945 3785 9975 3790
rect 9945 3765 9950 3785
rect 9970 3765 9975 3785
rect 9945 3760 9975 3765
rect 9950 3755 9970 3760
rect 10040 3625 10060 4080
rect 10085 3950 10105 4215
rect 10130 4195 10150 4200
rect 10125 4190 10155 4195
rect 10125 4170 10130 4190
rect 10150 4170 10155 4190
rect 10125 4165 10155 4170
rect 10080 3945 10110 3950
rect 10080 3925 10085 3945
rect 10105 3925 10110 3945
rect 10080 3920 10110 3925
rect 10085 3915 10105 3920
rect 10130 3910 10150 4165
rect 10175 3910 10195 4215
rect 10265 3950 10285 4215
rect 10310 4195 10330 4200
rect 10305 4190 10335 4195
rect 10305 4170 10310 4190
rect 10330 4170 10335 4190
rect 10305 4165 10335 4170
rect 10260 3945 10290 3950
rect 10260 3925 10265 3945
rect 10285 3925 10290 3945
rect 10260 3920 10290 3925
rect 10265 3915 10285 3920
rect 10220 3910 10240 3915
rect 10310 3910 10330 4165
rect 10355 3910 10375 4215
rect 10445 3950 10465 4215
rect 10490 4195 10510 4200
rect 10670 4195 10690 4200
rect 10485 4190 10515 4195
rect 10485 4170 10490 4190
rect 10510 4170 10515 4190
rect 10485 4165 10515 4170
rect 10665 4190 10695 4195
rect 10665 4170 10670 4190
rect 10690 4170 10695 4190
rect 10665 4165 10695 4170
rect 10440 3945 10470 3950
rect 10440 3925 10445 3945
rect 10465 3925 10470 3945
rect 10440 3920 10470 3925
rect 10445 3915 10465 3920
rect 10400 3910 10420 3915
rect 10125 3905 10155 3910
rect 10125 3885 10130 3905
rect 10150 3885 10155 3905
rect 10125 3880 10155 3885
rect 10170 3905 10200 3910
rect 10170 3885 10175 3905
rect 10195 3885 10200 3905
rect 10170 3880 10200 3885
rect 10215 3905 10245 3910
rect 10215 3885 10220 3905
rect 10240 3885 10245 3905
rect 10215 3880 10245 3885
rect 10305 3905 10335 3910
rect 10305 3885 10310 3905
rect 10330 3885 10335 3905
rect 10305 3880 10335 3885
rect 10350 3905 10380 3910
rect 10350 3885 10355 3905
rect 10375 3885 10380 3905
rect 10350 3880 10380 3885
rect 10395 3905 10425 3910
rect 10395 3885 10400 3905
rect 10420 3885 10425 3905
rect 10395 3880 10425 3885
rect 10130 3875 10150 3880
rect 10085 3830 10105 3835
rect 10080 3825 10110 3830
rect 10080 3805 10085 3825
rect 10105 3805 10110 3825
rect 10080 3800 10110 3805
rect 10035 3620 10065 3625
rect 10035 3600 10040 3620
rect 10060 3600 10065 3620
rect 10035 3595 10065 3600
rect 10040 3590 10060 3595
rect 10085 3575 10105 3800
rect 10175 3575 10195 3880
rect 10220 3625 10240 3880
rect 10310 3875 10330 3880
rect 10265 3830 10285 3835
rect 10260 3825 10290 3830
rect 10260 3805 10265 3825
rect 10285 3805 10290 3825
rect 10260 3800 10290 3805
rect 10215 3620 10245 3625
rect 10215 3600 10220 3620
rect 10240 3600 10245 3620
rect 10215 3595 10245 3600
rect 10220 3590 10240 3595
rect 10265 3575 10285 3800
rect 10355 3575 10375 3880
rect 10400 3625 10420 3880
rect 10445 3830 10465 3835
rect 10440 3825 10470 3830
rect 10440 3805 10445 3825
rect 10465 3805 10470 3825
rect 10440 3800 10470 3805
rect 10395 3620 10425 3625
rect 10395 3600 10400 3620
rect 10420 3600 10425 3620
rect 10395 3595 10425 3600
rect 10400 3590 10420 3595
rect 10445 3575 10465 3800
rect 10490 3790 10510 4165
rect 10580 4110 10600 4115
rect 10575 4105 10605 4110
rect 10575 4085 10580 4105
rect 10600 4085 10605 4105
rect 10575 4080 10605 4085
rect 10485 3785 10515 3790
rect 10485 3765 10490 3785
rect 10510 3765 10515 3785
rect 10485 3760 10515 3765
rect 10490 3755 10510 3760
rect 10580 3625 10600 4080
rect 10670 3790 10690 4165
rect 10760 4110 10780 4115
rect 10755 4105 10785 4110
rect 10755 4085 10760 4105
rect 10780 4085 10785 4105
rect 10755 4080 10785 4085
rect 10665 3785 10695 3790
rect 10665 3765 10670 3785
rect 10690 3765 10695 3785
rect 10665 3760 10695 3765
rect 10670 3755 10690 3760
rect 10760 3625 10780 4080
rect 10805 3950 10825 4215
rect 10850 4195 10870 4200
rect 10845 4190 10875 4195
rect 10845 4170 10850 4190
rect 10870 4170 10875 4190
rect 10845 4165 10875 4170
rect 10800 3945 10830 3950
rect 10800 3925 10805 3945
rect 10825 3925 10830 3945
rect 10800 3920 10830 3925
rect 10805 3915 10825 3920
rect 10850 3910 10870 4165
rect 10895 3910 10915 4215
rect 10985 3950 11005 4215
rect 11030 4195 11050 4200
rect 11025 4190 11055 4195
rect 11025 4170 11030 4190
rect 11050 4170 11055 4190
rect 11025 4165 11055 4170
rect 10980 3945 11010 3950
rect 10980 3925 10985 3945
rect 11005 3925 11010 3945
rect 10980 3920 11010 3925
rect 10985 3915 11005 3920
rect 10940 3910 10960 3915
rect 11030 3910 11050 4165
rect 11075 3910 11095 4215
rect 11165 3950 11185 4215
rect 11210 4195 11230 4200
rect 11390 4195 11410 4200
rect 11205 4190 11235 4195
rect 11205 4170 11210 4190
rect 11230 4170 11235 4190
rect 11205 4165 11235 4170
rect 11385 4190 11415 4195
rect 11385 4170 11390 4190
rect 11410 4170 11415 4190
rect 11385 4165 11415 4170
rect 11160 3945 11190 3950
rect 11160 3925 11165 3945
rect 11185 3925 11190 3945
rect 11160 3920 11190 3925
rect 11165 3915 11185 3920
rect 11120 3910 11140 3915
rect 10845 3905 10875 3910
rect 10845 3885 10850 3905
rect 10870 3885 10875 3905
rect 10845 3880 10875 3885
rect 10890 3905 10920 3910
rect 10890 3885 10895 3905
rect 10915 3885 10920 3905
rect 10890 3880 10920 3885
rect 10935 3905 10965 3910
rect 10935 3885 10940 3905
rect 10960 3885 10965 3905
rect 10935 3880 10965 3885
rect 11025 3905 11055 3910
rect 11025 3885 11030 3905
rect 11050 3885 11055 3905
rect 11025 3880 11055 3885
rect 11070 3905 11100 3910
rect 11070 3885 11075 3905
rect 11095 3885 11100 3905
rect 11070 3880 11100 3885
rect 11115 3905 11145 3910
rect 11115 3885 11120 3905
rect 11140 3885 11145 3905
rect 11115 3880 11145 3885
rect 10850 3875 10870 3880
rect 10805 3830 10825 3835
rect 10800 3825 10830 3830
rect 10800 3805 10805 3825
rect 10825 3805 10830 3825
rect 10800 3800 10830 3805
rect 10575 3620 10605 3625
rect 10575 3600 10580 3620
rect 10600 3600 10605 3620
rect 10575 3595 10605 3600
rect 10755 3620 10785 3625
rect 10755 3600 10760 3620
rect 10780 3600 10785 3620
rect 10755 3595 10785 3600
rect 10580 3590 10600 3595
rect 10760 3590 10780 3595
rect 10805 3575 10825 3800
rect 10895 3575 10915 3880
rect 10940 3625 10960 3880
rect 11030 3875 11050 3880
rect 10985 3830 11005 3835
rect 10980 3825 11010 3830
rect 10980 3805 10985 3825
rect 11005 3805 11010 3825
rect 10980 3800 11010 3805
rect 10935 3620 10965 3625
rect 10935 3600 10940 3620
rect 10960 3600 10965 3620
rect 10935 3595 10965 3600
rect 10940 3590 10960 3595
rect 10985 3575 11005 3800
rect 11075 3575 11095 3880
rect 11120 3625 11140 3880
rect 11165 3830 11185 3835
rect 11160 3825 11190 3830
rect 11160 3805 11165 3825
rect 11185 3805 11190 3825
rect 11160 3800 11190 3805
rect 11115 3620 11145 3625
rect 11115 3600 11120 3620
rect 11140 3600 11145 3620
rect 11115 3595 11145 3600
rect 11120 3590 11140 3595
rect 11165 3575 11185 3800
rect 11210 3790 11230 4165
rect 11300 4110 11320 4115
rect 11295 4105 11325 4110
rect 11295 4085 11300 4105
rect 11320 4085 11325 4105
rect 11295 4080 11325 4085
rect 11205 3785 11235 3790
rect 11205 3765 11210 3785
rect 11230 3765 11235 3785
rect 11205 3760 11235 3765
rect 11210 3755 11230 3760
rect 11300 3625 11320 4080
rect 11390 3790 11410 4165
rect 11480 4110 11500 4115
rect 11475 4105 11505 4110
rect 11475 4085 11480 4105
rect 11500 4085 11505 4105
rect 11475 4080 11505 4085
rect 11385 3785 11415 3790
rect 11385 3765 11390 3785
rect 11410 3765 11415 3785
rect 11385 3760 11415 3765
rect 11390 3755 11410 3760
rect 11480 3625 11500 4080
rect 11525 3950 11545 4215
rect 11570 4195 11590 4200
rect 11565 4190 11595 4195
rect 11565 4170 11570 4190
rect 11590 4170 11595 4190
rect 11565 4165 11595 4170
rect 11520 3945 11550 3950
rect 11520 3925 11525 3945
rect 11545 3925 11550 3945
rect 11520 3920 11550 3925
rect 11525 3915 11545 3920
rect 11570 3910 11590 4165
rect 11615 3910 11635 4215
rect 11705 3950 11725 4215
rect 11750 4195 11770 4200
rect 11745 4190 11775 4195
rect 11745 4170 11750 4190
rect 11770 4170 11775 4190
rect 11745 4165 11775 4170
rect 11700 3945 11730 3950
rect 11700 3925 11705 3945
rect 11725 3925 11730 3945
rect 11700 3920 11730 3925
rect 11705 3915 11725 3920
rect 11660 3910 11680 3915
rect 11750 3910 11770 4165
rect 11795 3910 11815 4215
rect 11885 3950 11905 4215
rect 11930 4195 11950 4200
rect 12110 4195 12130 4200
rect 11925 4190 11955 4195
rect 11925 4170 11930 4190
rect 11950 4170 11955 4190
rect 11925 4165 11955 4170
rect 12105 4190 12135 4195
rect 12105 4170 12110 4190
rect 12130 4170 12135 4190
rect 12105 4165 12135 4170
rect 11880 3945 11910 3950
rect 11880 3925 11885 3945
rect 11905 3925 11910 3945
rect 11880 3920 11910 3925
rect 11885 3915 11905 3920
rect 11840 3910 11860 3915
rect 11565 3905 11595 3910
rect 11565 3885 11570 3905
rect 11590 3885 11595 3905
rect 11565 3880 11595 3885
rect 11610 3905 11640 3910
rect 11610 3885 11615 3905
rect 11635 3885 11640 3905
rect 11610 3880 11640 3885
rect 11655 3905 11685 3910
rect 11655 3885 11660 3905
rect 11680 3885 11685 3905
rect 11655 3880 11685 3885
rect 11745 3905 11775 3910
rect 11745 3885 11750 3905
rect 11770 3885 11775 3905
rect 11745 3880 11775 3885
rect 11790 3905 11820 3910
rect 11790 3885 11795 3905
rect 11815 3885 11820 3905
rect 11790 3880 11820 3885
rect 11835 3905 11865 3910
rect 11835 3885 11840 3905
rect 11860 3885 11865 3905
rect 11835 3880 11865 3885
rect 11570 3875 11590 3880
rect 11525 3830 11545 3835
rect 11520 3825 11550 3830
rect 11520 3805 11525 3825
rect 11545 3805 11550 3825
rect 11520 3800 11550 3805
rect 11295 3620 11325 3625
rect 11295 3600 11300 3620
rect 11320 3600 11325 3620
rect 11295 3595 11325 3600
rect 11475 3620 11505 3625
rect 11475 3600 11480 3620
rect 11500 3600 11505 3620
rect 11475 3595 11505 3600
rect 11300 3590 11320 3595
rect 11480 3590 11500 3595
rect 11525 3575 11545 3800
rect 11615 3575 11635 3880
rect 11660 3625 11680 3880
rect 11750 3875 11770 3880
rect 11705 3830 11725 3835
rect 11700 3825 11730 3830
rect 11700 3805 11705 3825
rect 11725 3805 11730 3825
rect 11700 3800 11730 3805
rect 11655 3620 11685 3625
rect 11655 3600 11660 3620
rect 11680 3600 11685 3620
rect 11655 3595 11685 3600
rect 11660 3590 11680 3595
rect 11705 3575 11725 3800
rect 11795 3575 11815 3880
rect 11840 3625 11860 3880
rect 11885 3830 11905 3835
rect 11880 3825 11910 3830
rect 11880 3805 11885 3825
rect 11905 3805 11910 3825
rect 11880 3800 11910 3805
rect 11835 3620 11865 3625
rect 11835 3600 11840 3620
rect 11860 3600 11865 3620
rect 11835 3595 11865 3600
rect 11840 3590 11860 3595
rect 11885 3575 11905 3800
rect 11930 3790 11950 4165
rect 12020 4110 12040 4115
rect 12015 4105 12045 4110
rect 12015 4085 12020 4105
rect 12040 4085 12045 4105
rect 12015 4080 12045 4085
rect 11925 3785 11955 3790
rect 11925 3765 11930 3785
rect 11950 3765 11955 3785
rect 11925 3760 11955 3765
rect 11930 3755 11950 3760
rect 12020 3625 12040 4080
rect 12110 3790 12130 4165
rect 12200 4110 12220 4115
rect 12195 4105 12225 4110
rect 12195 4085 12200 4105
rect 12220 4085 12225 4105
rect 12195 4080 12225 4085
rect 12105 3785 12135 3790
rect 12105 3765 12110 3785
rect 12130 3765 12135 3785
rect 12105 3760 12135 3765
rect 12110 3755 12130 3760
rect 12200 3625 12220 4080
rect 12245 3950 12265 4215
rect 12290 4195 12310 4200
rect 12285 4190 12315 4195
rect 12285 4170 12290 4190
rect 12310 4170 12315 4190
rect 12285 4165 12315 4170
rect 12240 3945 12270 3950
rect 12240 3925 12245 3945
rect 12265 3925 12270 3945
rect 12240 3920 12270 3925
rect 12245 3915 12265 3920
rect 12290 3910 12310 4165
rect 12335 3910 12355 4215
rect 12425 3950 12445 4215
rect 12470 4195 12490 4200
rect 12465 4190 12495 4195
rect 12465 4170 12470 4190
rect 12490 4170 12495 4190
rect 12465 4165 12495 4170
rect 12420 3945 12450 3950
rect 12420 3925 12425 3945
rect 12445 3925 12450 3945
rect 12420 3920 12450 3925
rect 12425 3915 12445 3920
rect 12380 3910 12400 3915
rect 12470 3910 12490 4165
rect 12515 3910 12535 4215
rect 12605 3950 12625 4215
rect 12650 4195 12670 4200
rect 12830 4195 12850 4200
rect 12645 4190 12675 4195
rect 12645 4170 12650 4190
rect 12670 4170 12675 4190
rect 12645 4165 12675 4170
rect 12825 4190 12855 4195
rect 12825 4170 12830 4190
rect 12850 4170 12855 4190
rect 12825 4165 12855 4170
rect 12600 3945 12630 3950
rect 12600 3925 12605 3945
rect 12625 3925 12630 3945
rect 12600 3920 12630 3925
rect 12605 3915 12625 3920
rect 12560 3910 12580 3915
rect 12285 3905 12315 3910
rect 12285 3885 12290 3905
rect 12310 3885 12315 3905
rect 12285 3880 12315 3885
rect 12330 3905 12360 3910
rect 12330 3885 12335 3905
rect 12355 3885 12360 3905
rect 12330 3880 12360 3885
rect 12375 3905 12405 3910
rect 12375 3885 12380 3905
rect 12400 3885 12405 3905
rect 12375 3880 12405 3885
rect 12465 3905 12495 3910
rect 12465 3885 12470 3905
rect 12490 3885 12495 3905
rect 12465 3880 12495 3885
rect 12510 3905 12540 3910
rect 12510 3885 12515 3905
rect 12535 3885 12540 3905
rect 12510 3880 12540 3885
rect 12555 3905 12585 3910
rect 12555 3885 12560 3905
rect 12580 3885 12585 3905
rect 12555 3880 12585 3885
rect 12290 3875 12310 3880
rect 12245 3830 12265 3835
rect 12240 3825 12270 3830
rect 12240 3805 12245 3825
rect 12265 3805 12270 3825
rect 12240 3800 12270 3805
rect 12015 3620 12045 3625
rect 12015 3600 12020 3620
rect 12040 3600 12045 3620
rect 12015 3595 12045 3600
rect 12195 3620 12225 3625
rect 12195 3600 12200 3620
rect 12220 3600 12225 3620
rect 12195 3595 12225 3600
rect 12020 3590 12040 3595
rect 12200 3590 12220 3595
rect 12245 3575 12265 3800
rect 12335 3575 12355 3880
rect 12380 3625 12400 3880
rect 12470 3875 12490 3880
rect 12425 3830 12445 3835
rect 12420 3825 12450 3830
rect 12420 3805 12425 3825
rect 12445 3805 12450 3825
rect 12420 3800 12450 3805
rect 12375 3620 12405 3625
rect 12375 3600 12380 3620
rect 12400 3600 12405 3620
rect 12375 3595 12405 3600
rect 12380 3590 12400 3595
rect 12425 3575 12445 3800
rect 12515 3575 12535 3880
rect 12560 3625 12580 3880
rect 12605 3830 12625 3835
rect 12600 3825 12630 3830
rect 12600 3805 12605 3825
rect 12625 3805 12630 3825
rect 12600 3800 12630 3805
rect 12555 3620 12585 3625
rect 12555 3600 12560 3620
rect 12580 3600 12585 3620
rect 12555 3595 12585 3600
rect 12560 3590 12580 3595
rect 12605 3575 12625 3800
rect 12650 3790 12670 4165
rect 12740 4110 12760 4115
rect 12735 4105 12765 4110
rect 12735 4085 12740 4105
rect 12760 4085 12765 4105
rect 12735 4080 12765 4085
rect 12645 3785 12675 3790
rect 12645 3765 12650 3785
rect 12670 3765 12675 3785
rect 12645 3760 12675 3765
rect 12650 3755 12670 3760
rect 12740 3625 12760 4080
rect 12830 3790 12850 4165
rect 12920 4110 12940 4115
rect 12915 4105 12945 4110
rect 12915 4085 12920 4105
rect 12940 4085 12945 4105
rect 12915 4080 12945 4085
rect 12825 3785 12855 3790
rect 12825 3765 12830 3785
rect 12850 3765 12855 3785
rect 12825 3760 12855 3765
rect 12830 3755 12850 3760
rect 12920 3625 12940 4080
rect 12965 3950 12985 4215
rect 13010 4195 13030 4200
rect 13005 4190 13035 4195
rect 13005 4170 13010 4190
rect 13030 4170 13035 4190
rect 13005 4165 13035 4170
rect 12960 3945 12990 3950
rect 12960 3925 12965 3945
rect 12985 3925 12990 3945
rect 12960 3920 12990 3925
rect 12965 3915 12985 3920
rect 13010 3910 13030 4165
rect 13055 3910 13075 4215
rect 13145 3950 13165 4215
rect 13190 4195 13210 4200
rect 13185 4190 13215 4195
rect 13185 4170 13190 4190
rect 13210 4170 13215 4190
rect 13185 4165 13215 4170
rect 13140 3945 13170 3950
rect 13140 3925 13145 3945
rect 13165 3925 13170 3945
rect 13140 3920 13170 3925
rect 13145 3915 13165 3920
rect 13100 3910 13120 3915
rect 13190 3910 13210 4165
rect 13235 3910 13255 4215
rect 13325 3950 13345 4215
rect 13685 4210 13705 4215
rect 13370 4195 13390 4200
rect 13550 4195 13570 4200
rect 13730 4195 13750 4200
rect 13365 4190 13395 4195
rect 13365 4170 13370 4190
rect 13390 4170 13395 4190
rect 13365 4165 13395 4170
rect 13545 4190 13575 4195
rect 13545 4170 13550 4190
rect 13570 4170 13575 4190
rect 13545 4165 13575 4170
rect 13725 4190 13755 4195
rect 13725 4170 13730 4190
rect 13750 4170 13755 4190
rect 13725 4165 13755 4170
rect 13320 3945 13350 3950
rect 13320 3925 13325 3945
rect 13345 3925 13350 3945
rect 13320 3920 13350 3925
rect 13325 3915 13345 3920
rect 13280 3910 13300 3915
rect 13005 3905 13035 3910
rect 13005 3885 13010 3905
rect 13030 3885 13035 3905
rect 13005 3880 13035 3885
rect 13050 3905 13080 3910
rect 13050 3885 13055 3905
rect 13075 3885 13080 3905
rect 13050 3880 13080 3885
rect 13095 3905 13125 3910
rect 13095 3885 13100 3905
rect 13120 3885 13125 3905
rect 13095 3880 13125 3885
rect 13185 3905 13215 3910
rect 13185 3885 13190 3905
rect 13210 3885 13215 3905
rect 13185 3880 13215 3885
rect 13230 3905 13260 3910
rect 13230 3885 13235 3905
rect 13255 3885 13260 3905
rect 13230 3880 13260 3885
rect 13275 3905 13305 3910
rect 13275 3885 13280 3905
rect 13300 3885 13305 3905
rect 13275 3880 13305 3885
rect 13010 3875 13030 3880
rect 12965 3830 12985 3835
rect 12960 3825 12990 3830
rect 12960 3805 12965 3825
rect 12985 3805 12990 3825
rect 12960 3800 12990 3805
rect 12735 3620 12765 3625
rect 12735 3600 12740 3620
rect 12760 3600 12765 3620
rect 12735 3595 12765 3600
rect 12915 3620 12945 3625
rect 12915 3600 12920 3620
rect 12940 3600 12945 3620
rect 12915 3595 12945 3600
rect 12740 3590 12760 3595
rect 12920 3590 12940 3595
rect 12965 3575 12985 3800
rect 13055 3575 13075 3880
rect 13100 3625 13120 3880
rect 13190 3875 13210 3880
rect 13145 3830 13165 3835
rect 13140 3825 13170 3830
rect 13140 3805 13145 3825
rect 13165 3805 13170 3825
rect 13140 3800 13170 3805
rect 13095 3620 13125 3625
rect 13095 3600 13100 3620
rect 13120 3600 13125 3620
rect 13095 3595 13125 3600
rect 13100 3590 13120 3595
rect 13145 3575 13165 3800
rect 13235 3575 13255 3880
rect 13280 3625 13300 3880
rect 13325 3830 13345 3835
rect 13320 3825 13350 3830
rect 13320 3805 13325 3825
rect 13345 3805 13350 3825
rect 13320 3800 13350 3805
rect 13275 3620 13305 3625
rect 13275 3600 13280 3620
rect 13300 3600 13305 3620
rect 13275 3595 13305 3600
rect 13280 3590 13300 3595
rect 13325 3575 13345 3800
rect 13370 3790 13390 4165
rect 13460 4110 13480 4115
rect 13455 4105 13485 4110
rect 13455 4085 13460 4105
rect 13480 4085 13485 4105
rect 13455 4080 13485 4085
rect 13365 3785 13395 3790
rect 13365 3765 13370 3785
rect 13390 3765 13395 3785
rect 13365 3760 13395 3765
rect 13370 3755 13390 3760
rect 13460 3625 13480 4080
rect 13550 4030 13570 4165
rect 13640 4110 13660 4115
rect 13635 4105 13665 4110
rect 13635 4085 13640 4105
rect 13660 4085 13665 4105
rect 13635 4080 13665 4085
rect 13545 4025 13575 4030
rect 13545 4005 13550 4025
rect 13570 4005 13575 4025
rect 13545 4000 13575 4005
rect 13550 3995 13570 4000
rect 13640 3625 13660 4080
rect 13730 3990 13750 4165
rect 13775 4110 13795 4115
rect 13865 4110 13885 4215
rect 13910 4195 13930 4200
rect 14090 4195 14110 4200
rect 14270 4195 14290 4200
rect 13905 4190 13935 4195
rect 13905 4170 13910 4190
rect 13930 4170 13935 4190
rect 13905 4165 13935 4170
rect 14085 4190 14115 4195
rect 14085 4170 14090 4190
rect 14110 4170 14115 4190
rect 14085 4165 14115 4170
rect 14265 4190 14295 4195
rect 14265 4170 14270 4190
rect 14290 4170 14295 4190
rect 14265 4165 14295 4170
rect 13770 4105 13800 4110
rect 13770 4085 13775 4105
rect 13795 4085 13800 4105
rect 13770 4080 13800 4085
rect 13860 4105 13890 4110
rect 13860 4085 13865 4105
rect 13885 4085 13890 4105
rect 13860 4080 13890 4085
rect 13725 3985 13755 3990
rect 13725 3965 13730 3985
rect 13750 3965 13755 3985
rect 13725 3960 13755 3965
rect 13730 3955 13750 3960
rect 13685 3830 13705 3835
rect 13680 3825 13710 3830
rect 13680 3805 13685 3825
rect 13705 3805 13710 3825
rect 13680 3800 13710 3805
rect 13455 3620 13485 3625
rect 13455 3600 13460 3620
rect 13480 3600 13485 3620
rect 13455 3595 13485 3600
rect 13635 3620 13665 3625
rect 13635 3600 13640 3620
rect 13660 3600 13665 3620
rect 13635 3595 13665 3600
rect 13460 3590 13480 3595
rect 13640 3590 13660 3595
rect 13685 3575 13705 3800
rect 13775 3575 13795 4080
rect 13865 4075 13885 4080
rect 13910 3990 13930 4165
rect 13955 4110 13975 4115
rect 13950 4105 13980 4110
rect 13950 4085 13955 4105
rect 13975 4085 13980 4105
rect 13950 4080 13980 4085
rect 13905 3985 13935 3990
rect 13905 3965 13910 3985
rect 13930 3965 13935 3985
rect 13905 3960 13935 3965
rect 13910 3955 13930 3960
rect 13820 3870 13840 3875
rect 13815 3865 13845 3870
rect 13815 3845 13820 3865
rect 13840 3845 13845 3865
rect 13815 3840 13845 3845
rect 13820 3625 13840 3840
rect 13865 3830 13885 3835
rect 13860 3825 13890 3830
rect 13860 3805 13865 3825
rect 13885 3805 13890 3825
rect 13860 3800 13890 3805
rect 13815 3620 13845 3625
rect 13815 3600 13820 3620
rect 13840 3600 13845 3620
rect 13815 3595 13845 3600
rect 13820 3590 13840 3595
rect 13865 3575 13885 3800
rect 13955 3575 13975 4080
rect 14090 4030 14110 4165
rect 14180 4110 14200 4115
rect 14175 4105 14205 4110
rect 14175 4085 14180 4105
rect 14200 4085 14205 4105
rect 14175 4080 14205 4085
rect 14085 4025 14115 4030
rect 14085 4005 14090 4025
rect 14110 4005 14115 4025
rect 14085 4000 14115 4005
rect 14090 3995 14110 4000
rect 14000 3870 14020 3875
rect 13995 3865 14025 3870
rect 13995 3845 14000 3865
rect 14020 3845 14025 3865
rect 13995 3840 14025 3845
rect 14000 3625 14020 3840
rect 14045 3830 14065 3835
rect 14040 3825 14070 3830
rect 14040 3805 14045 3825
rect 14065 3805 14070 3825
rect 14040 3800 14070 3805
rect 13995 3620 14025 3625
rect 13995 3600 14000 3620
rect 14020 3600 14025 3620
rect 13995 3595 14025 3600
rect 14000 3590 14020 3595
rect 14045 3575 14065 3800
rect 14180 3625 14200 4080
rect 14270 3790 14290 4165
rect 14405 3950 14425 4215
rect 14450 4195 14470 4200
rect 14445 4190 14475 4195
rect 14445 4170 14450 4190
rect 14470 4170 14475 4190
rect 14445 4165 14475 4170
rect 14400 3945 14430 3950
rect 14400 3925 14405 3945
rect 14425 3925 14430 3945
rect 14400 3920 14430 3925
rect 14405 3915 14425 3920
rect 14450 3870 14470 4165
rect 14445 3865 14475 3870
rect 14445 3845 14450 3865
rect 14470 3845 14475 3865
rect 14445 3840 14475 3845
rect 14450 3835 14470 3840
rect 14495 3790 14515 4215
rect 14585 3950 14605 4215
rect 14630 4195 14650 4200
rect 14625 4190 14655 4195
rect 14625 4170 14630 4190
rect 14650 4170 14655 4190
rect 14625 4165 14655 4170
rect 14580 3945 14610 3950
rect 14580 3925 14585 3945
rect 14605 3925 14610 3945
rect 14580 3920 14610 3925
rect 14585 3915 14605 3920
rect 14630 3870 14650 4165
rect 14625 3865 14655 3870
rect 14625 3845 14630 3865
rect 14650 3845 14655 3865
rect 14625 3840 14655 3845
rect 14630 3835 14650 3840
rect 14585 3790 14605 3795
rect 14675 3790 14695 4215
rect 14765 3950 14785 4215
rect 14810 4195 14830 4200
rect 15080 4195 15100 4200
rect 14805 4190 14835 4195
rect 14805 4170 14810 4190
rect 14830 4170 14835 4190
rect 14805 4165 14835 4170
rect 15075 4190 15105 4195
rect 15075 4170 15080 4190
rect 15100 4170 15105 4190
rect 15075 4165 15105 4170
rect 14760 3945 14790 3950
rect 14760 3925 14765 3945
rect 14785 3925 14790 3945
rect 14760 3920 14790 3925
rect 14765 3915 14785 3920
rect 14810 3790 14830 4165
rect 15080 3790 15100 4165
rect 15125 3950 15145 4215
rect 15120 3945 15150 3950
rect 15120 3925 15125 3945
rect 15145 3925 15150 3945
rect 15120 3920 15150 3925
rect 15125 3915 15145 3920
rect 15215 3790 15235 4215
rect 15260 4195 15280 4200
rect 15255 4190 15285 4195
rect 15255 4170 15260 4190
rect 15280 4170 15285 4190
rect 15255 4165 15285 4170
rect 15260 3870 15280 4165
rect 15305 3950 15325 4215
rect 15300 3945 15330 3950
rect 15300 3925 15305 3945
rect 15325 3925 15330 3945
rect 15300 3920 15330 3925
rect 15305 3915 15325 3920
rect 15255 3865 15285 3870
rect 15255 3845 15260 3865
rect 15280 3845 15285 3865
rect 15255 3840 15285 3845
rect 15260 3835 15280 3840
rect 15305 3790 15325 3795
rect 15395 3790 15415 4215
rect 15440 4195 15460 4200
rect 15435 4190 15465 4195
rect 15435 4170 15440 4190
rect 15460 4170 15465 4190
rect 15435 4165 15465 4170
rect 15440 3870 15460 4165
rect 15485 3950 15505 4215
rect 15620 4195 15640 4200
rect 15800 4195 15820 4200
rect 15980 4195 16000 4200
rect 15615 4190 15645 4195
rect 15615 4170 15620 4190
rect 15640 4170 15645 4190
rect 15615 4165 15645 4170
rect 15795 4190 15825 4195
rect 15795 4170 15800 4190
rect 15820 4170 15825 4190
rect 15795 4165 15825 4170
rect 15975 4190 16005 4195
rect 15975 4170 15980 4190
rect 16000 4170 16005 4190
rect 15975 4165 16005 4170
rect 15480 3945 15510 3950
rect 15480 3925 15485 3945
rect 15505 3925 15510 3945
rect 15480 3920 15510 3925
rect 15485 3915 15505 3920
rect 15435 3865 15465 3870
rect 15435 3845 15440 3865
rect 15460 3845 15465 3865
rect 15435 3840 15465 3845
rect 15440 3835 15460 3840
rect 15620 3790 15640 4165
rect 15710 4110 15730 4115
rect 15705 4105 15735 4110
rect 15705 4085 15710 4105
rect 15730 4085 15735 4105
rect 15705 4080 15735 4085
rect 14265 3785 14295 3790
rect 14265 3765 14270 3785
rect 14290 3765 14295 3785
rect 14265 3760 14295 3765
rect 14490 3785 14520 3790
rect 14490 3765 14495 3785
rect 14515 3765 14520 3785
rect 14490 3760 14520 3765
rect 14580 3785 14610 3790
rect 14580 3765 14585 3785
rect 14605 3765 14610 3785
rect 14580 3760 14610 3765
rect 14670 3785 14700 3790
rect 14670 3765 14675 3785
rect 14695 3765 14700 3785
rect 14670 3760 14700 3765
rect 14805 3785 14835 3790
rect 14805 3765 14810 3785
rect 14830 3765 14835 3785
rect 14805 3760 14835 3765
rect 15075 3785 15105 3790
rect 15075 3765 15080 3785
rect 15100 3765 15105 3785
rect 15075 3760 15105 3765
rect 15210 3785 15240 3790
rect 15210 3765 15215 3785
rect 15235 3765 15240 3785
rect 15210 3760 15240 3765
rect 15300 3785 15330 3790
rect 15300 3765 15305 3785
rect 15325 3765 15330 3785
rect 15300 3760 15330 3765
rect 15390 3785 15420 3790
rect 15390 3765 15395 3785
rect 15415 3765 15420 3785
rect 15390 3760 15420 3765
rect 15615 3785 15645 3790
rect 15615 3765 15620 3785
rect 15640 3765 15645 3785
rect 15615 3760 15645 3765
rect 14270 3755 14290 3760
rect 14495 3755 14515 3760
rect 14540 3750 14560 3755
rect 14535 3745 14565 3750
rect 14535 3725 14540 3745
rect 14560 3725 14565 3745
rect 14535 3720 14565 3725
rect 14360 3710 14380 3715
rect 14355 3705 14385 3710
rect 14355 3685 14360 3705
rect 14380 3685 14385 3705
rect 14355 3680 14385 3685
rect 14360 3625 14380 3680
rect 14540 3625 14560 3720
rect 14175 3620 14205 3625
rect 14175 3600 14180 3620
rect 14200 3600 14205 3620
rect 14175 3595 14205 3600
rect 14355 3620 14385 3625
rect 14355 3600 14360 3620
rect 14380 3600 14385 3620
rect 14355 3595 14385 3600
rect 14535 3620 14565 3625
rect 14535 3600 14540 3620
rect 14560 3600 14565 3620
rect 14535 3595 14565 3600
rect 14180 3590 14200 3595
rect 14360 3590 14380 3595
rect 14540 3590 14560 3595
rect 14585 3575 14605 3760
rect 14675 3755 14695 3760
rect 14810 3755 14830 3760
rect 15080 3755 15100 3760
rect 15215 3755 15235 3760
rect 14720 3750 14740 3755
rect 15170 3750 15190 3755
rect 14715 3745 14745 3750
rect 14715 3725 14720 3745
rect 14740 3725 14745 3745
rect 14715 3720 14745 3725
rect 15165 3745 15195 3750
rect 15165 3725 15170 3745
rect 15190 3725 15195 3745
rect 15165 3720 15195 3725
rect 14720 3625 14740 3720
rect 14900 3710 14920 3715
rect 14990 3710 15010 3715
rect 14895 3705 14925 3710
rect 14895 3685 14900 3705
rect 14920 3685 14925 3705
rect 14895 3680 14925 3685
rect 14985 3705 15015 3710
rect 14985 3685 14990 3705
rect 15010 3685 15015 3705
rect 14985 3680 15015 3685
rect 14900 3625 14920 3680
rect 14990 3625 15010 3680
rect 15170 3625 15190 3720
rect 14715 3620 14745 3625
rect 14715 3600 14720 3620
rect 14740 3600 14745 3620
rect 14715 3595 14745 3600
rect 14895 3620 14925 3625
rect 14895 3600 14900 3620
rect 14920 3600 14925 3620
rect 14895 3595 14925 3600
rect 14985 3620 15015 3625
rect 14985 3600 14990 3620
rect 15010 3600 15015 3620
rect 14985 3595 15015 3600
rect 15165 3620 15195 3625
rect 15165 3600 15170 3620
rect 15190 3600 15195 3620
rect 15165 3595 15195 3600
rect 14720 3590 14740 3595
rect 14900 3590 14920 3595
rect 14990 3590 15010 3595
rect 15170 3590 15190 3595
rect 15305 3575 15325 3760
rect 15395 3755 15415 3760
rect 15620 3755 15640 3760
rect 15350 3750 15370 3755
rect 15345 3745 15375 3750
rect 15345 3725 15350 3745
rect 15370 3725 15375 3745
rect 15345 3720 15375 3725
rect 15350 3625 15370 3720
rect 15530 3710 15550 3715
rect 15525 3705 15555 3710
rect 15525 3685 15530 3705
rect 15550 3685 15555 3705
rect 15525 3680 15555 3685
rect 15530 3625 15550 3680
rect 15710 3625 15730 4080
rect 15800 4030 15820 4165
rect 15935 4110 15955 4115
rect 15930 4105 15960 4110
rect 15930 4085 15935 4105
rect 15955 4085 15960 4105
rect 15930 4080 15960 4085
rect 15795 4025 15825 4030
rect 15795 4005 15800 4025
rect 15820 4005 15825 4025
rect 15795 4000 15825 4005
rect 15800 3995 15820 4000
rect 15890 3870 15910 3875
rect 15885 3865 15915 3870
rect 15885 3845 15890 3865
rect 15910 3845 15915 3865
rect 15885 3840 15915 3845
rect 15845 3830 15865 3835
rect 15840 3825 15870 3830
rect 15840 3805 15845 3825
rect 15865 3805 15870 3825
rect 15840 3800 15870 3805
rect 15345 3620 15375 3625
rect 15345 3600 15350 3620
rect 15370 3600 15375 3620
rect 15345 3595 15375 3600
rect 15525 3620 15555 3625
rect 15525 3600 15530 3620
rect 15550 3600 15555 3620
rect 15525 3595 15555 3600
rect 15705 3620 15735 3625
rect 15705 3600 15710 3620
rect 15730 3600 15735 3620
rect 15705 3595 15735 3600
rect 15350 3590 15370 3595
rect 15530 3590 15550 3595
rect 15710 3590 15730 3595
rect 15845 3575 15865 3800
rect 15890 3625 15910 3840
rect 15885 3620 15915 3625
rect 15885 3600 15890 3620
rect 15910 3600 15915 3620
rect 15885 3595 15915 3600
rect 15890 3590 15910 3595
rect 15935 3575 15955 4080
rect 15980 3990 16000 4165
rect 16025 4110 16045 4215
rect 16205 4210 16225 4215
rect 16160 4195 16180 4200
rect 16340 4195 16360 4200
rect 16520 4195 16540 4200
rect 16155 4190 16185 4195
rect 16155 4170 16160 4190
rect 16180 4170 16185 4190
rect 16155 4165 16185 4170
rect 16335 4190 16365 4195
rect 16335 4170 16340 4190
rect 16360 4170 16365 4190
rect 16335 4165 16365 4170
rect 16515 4190 16545 4195
rect 16515 4170 16520 4190
rect 16540 4170 16545 4190
rect 16515 4165 16545 4170
rect 16115 4110 16135 4115
rect 16020 4105 16050 4110
rect 16020 4085 16025 4105
rect 16045 4085 16050 4105
rect 16020 4080 16050 4085
rect 16110 4105 16140 4110
rect 16110 4085 16115 4105
rect 16135 4085 16140 4105
rect 16110 4080 16140 4085
rect 16025 4075 16045 4080
rect 15975 3985 16005 3990
rect 15975 3965 15980 3985
rect 16000 3965 16005 3985
rect 15975 3960 16005 3965
rect 15980 3955 16000 3960
rect 16070 3870 16090 3875
rect 16065 3865 16095 3870
rect 16065 3845 16070 3865
rect 16090 3845 16095 3865
rect 16065 3840 16095 3845
rect 16025 3830 16045 3835
rect 16020 3825 16050 3830
rect 16020 3805 16025 3825
rect 16045 3805 16050 3825
rect 16020 3800 16050 3805
rect 16025 3575 16045 3800
rect 16070 3625 16090 3840
rect 16065 3620 16095 3625
rect 16065 3600 16070 3620
rect 16090 3600 16095 3620
rect 16065 3595 16095 3600
rect 16070 3590 16090 3595
rect 16115 3575 16135 4080
rect 16160 3990 16180 4165
rect 16250 4110 16270 4115
rect 16245 4105 16275 4110
rect 16245 4085 16250 4105
rect 16270 4085 16275 4105
rect 16245 4080 16275 4085
rect 16155 3985 16185 3990
rect 16155 3965 16160 3985
rect 16180 3965 16185 3985
rect 16155 3960 16185 3965
rect 16160 3955 16180 3960
rect 16205 3830 16225 3835
rect 16200 3825 16230 3830
rect 16200 3805 16205 3825
rect 16225 3805 16230 3825
rect 16200 3800 16230 3805
rect 16205 3575 16225 3800
rect 16250 3625 16270 4080
rect 16340 4030 16360 4165
rect 16430 4110 16450 4115
rect 16425 4105 16455 4110
rect 16425 4085 16430 4105
rect 16450 4085 16455 4105
rect 16425 4080 16455 4085
rect 16335 4025 16365 4030
rect 16335 4005 16340 4025
rect 16360 4005 16365 4025
rect 16335 4000 16365 4005
rect 16340 3995 16360 4000
rect 16430 3625 16450 4080
rect 16520 3790 16540 4165
rect 16565 3950 16585 4215
rect 16560 3945 16590 3950
rect 16560 3925 16565 3945
rect 16585 3925 16590 3945
rect 16560 3920 16590 3925
rect 16565 3915 16585 3920
rect 16610 3910 16630 3915
rect 16655 3910 16675 4215
rect 16700 4195 16720 4200
rect 16695 4190 16725 4195
rect 16695 4170 16700 4190
rect 16720 4170 16725 4190
rect 16695 4165 16725 4170
rect 16700 3910 16720 4165
rect 16745 3950 16765 4215
rect 16740 3945 16770 3950
rect 16740 3925 16745 3945
rect 16765 3925 16770 3945
rect 16740 3920 16770 3925
rect 16745 3915 16765 3920
rect 16790 3910 16810 3915
rect 16835 3910 16855 4215
rect 16880 4195 16900 4200
rect 16875 4190 16905 4195
rect 16875 4170 16880 4190
rect 16900 4170 16905 4190
rect 16875 4165 16905 4170
rect 16880 3910 16900 4165
rect 16925 3950 16945 4215
rect 17060 4195 17080 4200
rect 17240 4195 17260 4200
rect 17055 4190 17085 4195
rect 17055 4170 17060 4190
rect 17080 4170 17085 4190
rect 17055 4165 17085 4170
rect 17235 4190 17265 4195
rect 17235 4170 17240 4190
rect 17260 4170 17265 4190
rect 17235 4165 17265 4170
rect 16970 4110 16990 4115
rect 16965 4105 16995 4110
rect 16965 4085 16970 4105
rect 16990 4085 16995 4105
rect 16965 4080 16995 4085
rect 16920 3945 16950 3950
rect 16920 3925 16925 3945
rect 16945 3925 16950 3945
rect 16920 3920 16950 3925
rect 16925 3915 16945 3920
rect 16605 3905 16635 3910
rect 16605 3885 16610 3905
rect 16630 3885 16635 3905
rect 16605 3880 16635 3885
rect 16650 3905 16680 3910
rect 16650 3885 16655 3905
rect 16675 3885 16680 3905
rect 16650 3880 16680 3885
rect 16695 3905 16725 3910
rect 16695 3885 16700 3905
rect 16720 3885 16725 3905
rect 16695 3880 16725 3885
rect 16785 3905 16815 3910
rect 16785 3885 16790 3905
rect 16810 3885 16815 3905
rect 16785 3880 16815 3885
rect 16830 3905 16860 3910
rect 16830 3885 16835 3905
rect 16855 3885 16860 3905
rect 16830 3880 16860 3885
rect 16875 3905 16905 3910
rect 16875 3885 16880 3905
rect 16900 3885 16905 3905
rect 16875 3880 16905 3885
rect 16565 3830 16585 3835
rect 16560 3825 16590 3830
rect 16560 3805 16565 3825
rect 16585 3805 16590 3825
rect 16560 3800 16590 3805
rect 16515 3785 16545 3790
rect 16515 3765 16520 3785
rect 16540 3765 16545 3785
rect 16515 3760 16545 3765
rect 16520 3755 16540 3760
rect 16245 3620 16275 3625
rect 16245 3600 16250 3620
rect 16270 3600 16275 3620
rect 16245 3595 16275 3600
rect 16425 3620 16455 3625
rect 16425 3600 16430 3620
rect 16450 3600 16455 3620
rect 16425 3595 16455 3600
rect 16250 3590 16270 3595
rect 16430 3590 16450 3595
rect 16565 3575 16585 3800
rect 16610 3625 16630 3880
rect 16605 3620 16635 3625
rect 16605 3600 16610 3620
rect 16630 3600 16635 3620
rect 16605 3595 16635 3600
rect 16610 3590 16630 3595
rect 16655 3575 16675 3880
rect 16700 3875 16720 3880
rect 16745 3830 16765 3835
rect 16740 3825 16770 3830
rect 16740 3805 16745 3825
rect 16765 3805 16770 3825
rect 16740 3800 16770 3805
rect 16745 3575 16765 3800
rect 16790 3625 16810 3880
rect 16785 3620 16815 3625
rect 16785 3600 16790 3620
rect 16810 3600 16815 3620
rect 16785 3595 16815 3600
rect 16790 3590 16810 3595
rect 16835 3575 16855 3880
rect 16880 3875 16900 3880
rect 16925 3830 16945 3835
rect 16920 3825 16950 3830
rect 16920 3805 16925 3825
rect 16945 3805 16950 3825
rect 16920 3800 16950 3805
rect 16925 3575 16945 3800
rect 16970 3625 16990 4080
rect 17060 3790 17080 4165
rect 17150 4110 17170 4115
rect 17145 4105 17175 4110
rect 17145 4085 17150 4105
rect 17170 4085 17175 4105
rect 17145 4080 17175 4085
rect 17055 3785 17085 3790
rect 17055 3765 17060 3785
rect 17080 3765 17085 3785
rect 17055 3760 17085 3765
rect 17060 3755 17080 3760
rect 17150 3625 17170 4080
rect 17240 3790 17260 4165
rect 17285 3950 17305 4215
rect 17280 3945 17310 3950
rect 17280 3925 17285 3945
rect 17305 3925 17310 3945
rect 17280 3920 17310 3925
rect 17285 3915 17305 3920
rect 17330 3910 17350 3915
rect 17375 3910 17395 4215
rect 17420 4195 17440 4200
rect 17415 4190 17445 4195
rect 17415 4170 17420 4190
rect 17440 4170 17445 4190
rect 17415 4165 17445 4170
rect 17420 3910 17440 4165
rect 17465 3950 17485 4215
rect 17460 3945 17490 3950
rect 17460 3925 17465 3945
rect 17485 3925 17490 3945
rect 17460 3920 17490 3925
rect 17465 3915 17485 3920
rect 17510 3910 17530 3915
rect 17555 3910 17575 4215
rect 17600 4195 17620 4200
rect 17595 4190 17625 4195
rect 17595 4170 17600 4190
rect 17620 4170 17625 4190
rect 17595 4165 17625 4170
rect 17600 3910 17620 4165
rect 17645 3950 17665 4215
rect 17780 4195 17800 4200
rect 17960 4195 17980 4200
rect 17775 4190 17805 4195
rect 17775 4170 17780 4190
rect 17800 4170 17805 4190
rect 17775 4165 17805 4170
rect 17955 4190 17985 4195
rect 17955 4170 17960 4190
rect 17980 4170 17985 4190
rect 17955 4165 17985 4170
rect 17690 4110 17710 4115
rect 17685 4105 17715 4110
rect 17685 4085 17690 4105
rect 17710 4085 17715 4105
rect 17685 4080 17715 4085
rect 17640 3945 17670 3950
rect 17640 3925 17645 3945
rect 17665 3925 17670 3945
rect 17640 3920 17670 3925
rect 17645 3915 17665 3920
rect 17325 3905 17355 3910
rect 17325 3885 17330 3905
rect 17350 3885 17355 3905
rect 17325 3880 17355 3885
rect 17370 3905 17400 3910
rect 17370 3885 17375 3905
rect 17395 3885 17400 3905
rect 17370 3880 17400 3885
rect 17415 3905 17445 3910
rect 17415 3885 17420 3905
rect 17440 3885 17445 3905
rect 17415 3880 17445 3885
rect 17505 3905 17535 3910
rect 17505 3885 17510 3905
rect 17530 3885 17535 3905
rect 17505 3880 17535 3885
rect 17550 3905 17580 3910
rect 17550 3885 17555 3905
rect 17575 3885 17580 3905
rect 17550 3880 17580 3885
rect 17595 3905 17625 3910
rect 17595 3885 17600 3905
rect 17620 3885 17625 3905
rect 17595 3880 17625 3885
rect 17285 3830 17305 3835
rect 17280 3825 17310 3830
rect 17280 3805 17285 3825
rect 17305 3805 17310 3825
rect 17280 3800 17310 3805
rect 17235 3785 17265 3790
rect 17235 3765 17240 3785
rect 17260 3765 17265 3785
rect 17235 3760 17265 3765
rect 17240 3755 17260 3760
rect 16965 3620 16995 3625
rect 16965 3600 16970 3620
rect 16990 3600 16995 3620
rect 16965 3595 16995 3600
rect 17145 3620 17175 3625
rect 17145 3600 17150 3620
rect 17170 3600 17175 3620
rect 17145 3595 17175 3600
rect 16970 3590 16990 3595
rect 17150 3590 17170 3595
rect 17285 3575 17305 3800
rect 17330 3625 17350 3880
rect 17325 3620 17355 3625
rect 17325 3600 17330 3620
rect 17350 3600 17355 3620
rect 17325 3595 17355 3600
rect 17330 3590 17350 3595
rect 17375 3575 17395 3880
rect 17420 3875 17440 3880
rect 17465 3830 17485 3835
rect 17460 3825 17490 3830
rect 17460 3805 17465 3825
rect 17485 3805 17490 3825
rect 17460 3800 17490 3805
rect 17465 3575 17485 3800
rect 17510 3625 17530 3880
rect 17505 3620 17535 3625
rect 17505 3600 17510 3620
rect 17530 3600 17535 3620
rect 17505 3595 17535 3600
rect 17510 3590 17530 3595
rect 17555 3575 17575 3880
rect 17600 3875 17620 3880
rect 17645 3830 17665 3835
rect 17640 3825 17670 3830
rect 17640 3805 17645 3825
rect 17665 3805 17670 3825
rect 17640 3800 17670 3805
rect 17645 3575 17665 3800
rect 17690 3625 17710 4080
rect 17780 3790 17800 4165
rect 17870 4110 17890 4115
rect 17865 4105 17895 4110
rect 17865 4085 17870 4105
rect 17890 4085 17895 4105
rect 17865 4080 17895 4085
rect 17775 3785 17805 3790
rect 17775 3765 17780 3785
rect 17800 3765 17805 3785
rect 17775 3760 17805 3765
rect 17780 3755 17800 3760
rect 17870 3625 17890 4080
rect 17960 3790 17980 4165
rect 18005 3950 18025 4215
rect 18000 3945 18030 3950
rect 18000 3925 18005 3945
rect 18025 3925 18030 3945
rect 18000 3920 18030 3925
rect 18005 3915 18025 3920
rect 18050 3910 18070 3915
rect 18095 3910 18115 4215
rect 18140 4195 18160 4200
rect 18135 4190 18165 4195
rect 18135 4170 18140 4190
rect 18160 4170 18165 4190
rect 18135 4165 18165 4170
rect 18140 3910 18160 4165
rect 18185 3950 18205 4215
rect 18180 3945 18210 3950
rect 18180 3925 18185 3945
rect 18205 3925 18210 3945
rect 18180 3920 18210 3925
rect 18185 3915 18205 3920
rect 18230 3910 18250 3915
rect 18275 3910 18295 4215
rect 18320 4195 18340 4200
rect 18315 4190 18345 4195
rect 18315 4170 18320 4190
rect 18340 4170 18345 4190
rect 18315 4165 18345 4170
rect 18320 3910 18340 4165
rect 18365 3950 18385 4215
rect 18500 4195 18520 4200
rect 18680 4195 18700 4200
rect 18495 4190 18525 4195
rect 18495 4170 18500 4190
rect 18520 4170 18525 4190
rect 18495 4165 18525 4170
rect 18675 4190 18705 4195
rect 18675 4170 18680 4190
rect 18700 4170 18705 4190
rect 18675 4165 18705 4170
rect 18410 4110 18430 4115
rect 18405 4105 18435 4110
rect 18405 4085 18410 4105
rect 18430 4085 18435 4105
rect 18405 4080 18435 4085
rect 18360 3945 18390 3950
rect 18360 3925 18365 3945
rect 18385 3925 18390 3945
rect 18360 3920 18390 3925
rect 18365 3915 18385 3920
rect 18045 3905 18075 3910
rect 18045 3885 18050 3905
rect 18070 3885 18075 3905
rect 18045 3880 18075 3885
rect 18090 3905 18120 3910
rect 18090 3885 18095 3905
rect 18115 3885 18120 3905
rect 18090 3880 18120 3885
rect 18135 3905 18165 3910
rect 18135 3885 18140 3905
rect 18160 3885 18165 3905
rect 18135 3880 18165 3885
rect 18225 3905 18255 3910
rect 18225 3885 18230 3905
rect 18250 3885 18255 3905
rect 18225 3880 18255 3885
rect 18270 3905 18300 3910
rect 18270 3885 18275 3905
rect 18295 3885 18300 3905
rect 18270 3880 18300 3885
rect 18315 3905 18345 3910
rect 18315 3885 18320 3905
rect 18340 3885 18345 3905
rect 18315 3880 18345 3885
rect 18005 3830 18025 3835
rect 18000 3825 18030 3830
rect 18000 3805 18005 3825
rect 18025 3805 18030 3825
rect 18000 3800 18030 3805
rect 17955 3785 17985 3790
rect 17955 3765 17960 3785
rect 17980 3765 17985 3785
rect 17955 3760 17985 3765
rect 17960 3755 17980 3760
rect 17685 3620 17715 3625
rect 17685 3600 17690 3620
rect 17710 3600 17715 3620
rect 17685 3595 17715 3600
rect 17865 3620 17895 3625
rect 17865 3600 17870 3620
rect 17890 3600 17895 3620
rect 17865 3595 17895 3600
rect 17690 3590 17710 3595
rect 17870 3590 17890 3595
rect 18005 3575 18025 3800
rect 18050 3625 18070 3880
rect 18045 3620 18075 3625
rect 18045 3600 18050 3620
rect 18070 3600 18075 3620
rect 18045 3595 18075 3600
rect 18050 3590 18070 3595
rect 18095 3575 18115 3880
rect 18140 3875 18160 3880
rect 18185 3830 18205 3835
rect 18180 3825 18210 3830
rect 18180 3805 18185 3825
rect 18205 3805 18210 3825
rect 18180 3800 18210 3805
rect 18185 3575 18205 3800
rect 18230 3625 18250 3880
rect 18225 3620 18255 3625
rect 18225 3600 18230 3620
rect 18250 3600 18255 3620
rect 18225 3595 18255 3600
rect 18230 3590 18250 3595
rect 18275 3575 18295 3880
rect 18320 3875 18340 3880
rect 18365 3830 18385 3835
rect 18360 3825 18390 3830
rect 18360 3805 18365 3825
rect 18385 3805 18390 3825
rect 18360 3800 18390 3805
rect 18365 3575 18385 3800
rect 18410 3625 18430 4080
rect 18500 3790 18520 4165
rect 18590 4110 18610 4115
rect 18585 4105 18615 4110
rect 18585 4085 18590 4105
rect 18610 4085 18615 4105
rect 18585 4080 18615 4085
rect 18495 3785 18525 3790
rect 18495 3765 18500 3785
rect 18520 3765 18525 3785
rect 18495 3760 18525 3765
rect 18500 3755 18520 3760
rect 18590 3625 18610 4080
rect 18680 3790 18700 4165
rect 18725 3950 18745 4215
rect 18720 3945 18750 3950
rect 18720 3925 18725 3945
rect 18745 3925 18750 3945
rect 18720 3920 18750 3925
rect 18725 3915 18745 3920
rect 18770 3910 18790 3915
rect 18815 3910 18835 4215
rect 18860 4195 18880 4200
rect 18855 4190 18885 4195
rect 18855 4170 18860 4190
rect 18880 4170 18885 4190
rect 18855 4165 18885 4170
rect 18860 3910 18880 4165
rect 18905 3950 18925 4215
rect 18900 3945 18930 3950
rect 18900 3925 18905 3945
rect 18925 3925 18930 3945
rect 18900 3920 18930 3925
rect 18905 3915 18925 3920
rect 18950 3910 18970 3915
rect 18995 3910 19015 4215
rect 19040 4195 19060 4200
rect 19035 4190 19065 4195
rect 19035 4170 19040 4190
rect 19060 4170 19065 4190
rect 19035 4165 19065 4170
rect 19040 3910 19060 4165
rect 19085 3950 19105 4215
rect 19220 4195 19240 4200
rect 19400 4195 19420 4200
rect 19215 4190 19245 4195
rect 19215 4170 19220 4190
rect 19240 4170 19245 4190
rect 19215 4165 19245 4170
rect 19395 4190 19425 4195
rect 19395 4170 19400 4190
rect 19420 4170 19425 4190
rect 19395 4165 19425 4170
rect 19130 4110 19150 4115
rect 19125 4105 19155 4110
rect 19125 4085 19130 4105
rect 19150 4085 19155 4105
rect 19125 4080 19155 4085
rect 19080 3945 19110 3950
rect 19080 3925 19085 3945
rect 19105 3925 19110 3945
rect 19080 3920 19110 3925
rect 19085 3915 19105 3920
rect 18765 3905 18795 3910
rect 18765 3885 18770 3905
rect 18790 3885 18795 3905
rect 18765 3880 18795 3885
rect 18810 3905 18840 3910
rect 18810 3885 18815 3905
rect 18835 3885 18840 3905
rect 18810 3880 18840 3885
rect 18855 3905 18885 3910
rect 18855 3885 18860 3905
rect 18880 3885 18885 3905
rect 18855 3880 18885 3885
rect 18945 3905 18975 3910
rect 18945 3885 18950 3905
rect 18970 3885 18975 3905
rect 18945 3880 18975 3885
rect 18990 3905 19020 3910
rect 18990 3885 18995 3905
rect 19015 3885 19020 3905
rect 18990 3880 19020 3885
rect 19035 3905 19065 3910
rect 19035 3885 19040 3905
rect 19060 3885 19065 3905
rect 19035 3880 19065 3885
rect 18725 3830 18745 3835
rect 18720 3825 18750 3830
rect 18720 3805 18725 3825
rect 18745 3805 18750 3825
rect 18720 3800 18750 3805
rect 18675 3785 18705 3790
rect 18675 3765 18680 3785
rect 18700 3765 18705 3785
rect 18675 3760 18705 3765
rect 18680 3755 18700 3760
rect 18405 3620 18435 3625
rect 18405 3600 18410 3620
rect 18430 3600 18435 3620
rect 18405 3595 18435 3600
rect 18585 3620 18615 3625
rect 18585 3600 18590 3620
rect 18610 3600 18615 3620
rect 18585 3595 18615 3600
rect 18410 3590 18430 3595
rect 18590 3590 18610 3595
rect 18725 3575 18745 3800
rect 18770 3625 18790 3880
rect 18765 3620 18795 3625
rect 18765 3600 18770 3620
rect 18790 3600 18795 3620
rect 18765 3595 18795 3600
rect 18770 3590 18790 3595
rect 18815 3575 18835 3880
rect 18860 3875 18880 3880
rect 18905 3830 18925 3835
rect 18900 3825 18930 3830
rect 18900 3805 18905 3825
rect 18925 3805 18930 3825
rect 18900 3800 18930 3805
rect 18905 3575 18925 3800
rect 18950 3625 18970 3880
rect 18945 3620 18975 3625
rect 18945 3600 18950 3620
rect 18970 3600 18975 3620
rect 18945 3595 18975 3600
rect 18950 3590 18970 3595
rect 18995 3575 19015 3880
rect 19040 3875 19060 3880
rect 19085 3830 19105 3835
rect 19080 3825 19110 3830
rect 19080 3805 19085 3825
rect 19105 3805 19110 3825
rect 19080 3800 19110 3805
rect 19085 3575 19105 3800
rect 19130 3625 19150 4080
rect 19220 3790 19240 4165
rect 19310 4110 19330 4115
rect 19305 4105 19335 4110
rect 19305 4085 19310 4105
rect 19330 4085 19335 4105
rect 19305 4080 19335 4085
rect 19215 3785 19245 3790
rect 19215 3765 19220 3785
rect 19240 3765 19245 3785
rect 19215 3760 19245 3765
rect 19220 3755 19240 3760
rect 19310 3625 19330 4080
rect 19400 3790 19420 4165
rect 19445 3950 19465 4215
rect 19440 3945 19470 3950
rect 19440 3925 19445 3945
rect 19465 3925 19470 3945
rect 19440 3920 19470 3925
rect 19445 3915 19465 3920
rect 19490 3910 19510 3915
rect 19535 3910 19555 4215
rect 19580 4195 19600 4200
rect 19575 4190 19605 4195
rect 19575 4170 19580 4190
rect 19600 4170 19605 4190
rect 19575 4165 19605 4170
rect 19580 3910 19600 4165
rect 19625 3950 19645 4215
rect 19620 3945 19650 3950
rect 19620 3925 19625 3945
rect 19645 3925 19650 3945
rect 19620 3920 19650 3925
rect 19625 3915 19645 3920
rect 19670 3910 19690 3915
rect 19715 3910 19735 4215
rect 19760 4195 19780 4200
rect 19755 4190 19785 4195
rect 19755 4170 19760 4190
rect 19780 4170 19785 4190
rect 19755 4165 19785 4170
rect 19760 3910 19780 4165
rect 19805 3950 19825 4215
rect 19940 4195 19960 4200
rect 19935 4190 19965 4195
rect 19935 4170 19940 4190
rect 19960 4170 19965 4190
rect 19935 4165 19965 4170
rect 19850 4110 19870 4115
rect 19845 4105 19875 4110
rect 19845 4085 19850 4105
rect 19870 4085 19875 4105
rect 19845 4080 19875 4085
rect 19800 3945 19830 3950
rect 19800 3925 19805 3945
rect 19825 3925 19830 3945
rect 19800 3920 19830 3925
rect 19805 3915 19825 3920
rect 19485 3905 19515 3910
rect 19485 3885 19490 3905
rect 19510 3885 19515 3905
rect 19485 3880 19515 3885
rect 19530 3905 19560 3910
rect 19530 3885 19535 3905
rect 19555 3885 19560 3905
rect 19530 3880 19560 3885
rect 19575 3905 19605 3910
rect 19575 3885 19580 3905
rect 19600 3885 19605 3905
rect 19575 3880 19605 3885
rect 19665 3905 19695 3910
rect 19665 3885 19670 3905
rect 19690 3885 19695 3905
rect 19665 3880 19695 3885
rect 19710 3905 19740 3910
rect 19710 3885 19715 3905
rect 19735 3885 19740 3905
rect 19710 3880 19740 3885
rect 19755 3905 19785 3910
rect 19755 3885 19760 3905
rect 19780 3885 19785 3905
rect 19755 3880 19785 3885
rect 19445 3830 19465 3835
rect 19440 3825 19470 3830
rect 19440 3805 19445 3825
rect 19465 3805 19470 3825
rect 19440 3800 19470 3805
rect 19395 3785 19425 3790
rect 19395 3765 19400 3785
rect 19420 3765 19425 3785
rect 19395 3760 19425 3765
rect 19400 3755 19420 3760
rect 19125 3620 19155 3625
rect 19125 3600 19130 3620
rect 19150 3600 19155 3620
rect 19125 3595 19155 3600
rect 19305 3620 19335 3625
rect 19305 3600 19310 3620
rect 19330 3600 19335 3620
rect 19305 3595 19335 3600
rect 19130 3590 19150 3595
rect 19310 3590 19330 3595
rect 19445 3575 19465 3800
rect 19490 3625 19510 3880
rect 19485 3620 19515 3625
rect 19485 3600 19490 3620
rect 19510 3600 19515 3620
rect 19485 3595 19515 3600
rect 19490 3590 19510 3595
rect 19535 3575 19555 3880
rect 19580 3875 19600 3880
rect 19625 3830 19645 3835
rect 19620 3825 19650 3830
rect 19620 3805 19625 3825
rect 19645 3805 19650 3825
rect 19620 3800 19650 3805
rect 19625 3575 19645 3800
rect 19670 3625 19690 3880
rect 19665 3620 19695 3625
rect 19665 3600 19670 3620
rect 19690 3600 19695 3620
rect 19665 3595 19695 3600
rect 19670 3590 19690 3595
rect 19715 3575 19735 3880
rect 19760 3875 19780 3880
rect 19805 3830 19825 3835
rect 19800 3825 19830 3830
rect 19800 3805 19805 3825
rect 19825 3805 19830 3825
rect 19800 3800 19830 3805
rect 19805 3575 19825 3800
rect 19850 3625 19870 4080
rect 19940 3790 19960 4165
rect 19935 3785 19965 3790
rect 19935 3765 19940 3785
rect 19960 3765 19965 3785
rect 19935 3760 19965 3765
rect 19940 3755 19960 3760
rect 19845 3620 19875 3625
rect 19845 3600 19850 3620
rect 19870 3600 19875 3620
rect 19845 3595 19875 3600
rect 19850 3590 19870 3595
rect 20075 3575 20095 4215
rect 20165 3575 20185 4215
rect 20255 3575 20275 4215
rect 20345 4030 20365 4215
rect 20340 4025 20370 4030
rect 20340 4005 20345 4025
rect 20365 4005 20370 4025
rect 20340 4000 20370 4005
rect 20345 3575 20365 4000
rect 20435 3990 20455 4215
rect 20430 3985 20460 3990
rect 20430 3965 20435 3985
rect 20455 3965 20460 3985
rect 20430 3960 20460 3965
rect 20435 3575 20455 3960
rect 20525 3710 20545 4215
rect 20615 3750 20635 4215
rect 20610 3745 20640 3750
rect 20610 3725 20615 3745
rect 20635 3725 20640 3745
rect 20610 3720 20640 3725
rect 20520 3705 20550 3710
rect 20520 3685 20525 3705
rect 20545 3685 20550 3705
rect 20520 3680 20550 3685
rect 20525 3575 20545 3680
rect 20615 3575 20635 3720
rect 9180 3565 9210 3575
rect 9180 3485 9185 3565
rect 9205 3485 9210 3565
rect 9180 3475 9210 3485
rect 9270 3475 9300 3575
rect 9360 3475 9390 3575
rect 9450 3475 9480 3575
rect 9540 3475 9570 3575
rect 9630 3475 9660 3575
rect 9720 3475 9750 3575
rect 9810 3475 9840 3575
rect 9900 3565 9930 3575
rect 9900 3485 9905 3565
rect 9925 3485 9930 3565
rect 9900 3475 9930 3485
rect 9990 3565 10020 3575
rect 9990 3485 9995 3565
rect 10015 3485 10020 3565
rect 9990 3475 10020 3485
rect 10080 3565 10110 3575
rect 10080 3485 10085 3565
rect 10105 3485 10110 3565
rect 10080 3475 10110 3485
rect 10170 3565 10200 3575
rect 10170 3485 10175 3565
rect 10195 3485 10200 3565
rect 10170 3475 10200 3485
rect 10260 3565 10290 3575
rect 10260 3485 10265 3565
rect 10285 3485 10290 3565
rect 10260 3475 10290 3485
rect 10350 3565 10380 3575
rect 10350 3485 10355 3565
rect 10375 3485 10380 3565
rect 10350 3475 10380 3485
rect 10440 3565 10470 3575
rect 10440 3485 10445 3565
rect 10465 3485 10470 3565
rect 10440 3475 10470 3485
rect 10530 3565 10560 3575
rect 10530 3485 10535 3565
rect 10555 3485 10560 3565
rect 10530 3475 10560 3485
rect 10620 3565 10650 3575
rect 10620 3485 10625 3565
rect 10645 3485 10650 3565
rect 10620 3475 10650 3485
rect 10710 3565 10740 3575
rect 10710 3485 10715 3565
rect 10735 3485 10740 3565
rect 10710 3475 10740 3485
rect 10800 3565 10830 3575
rect 10800 3485 10805 3565
rect 10825 3485 10830 3565
rect 10800 3475 10830 3485
rect 10890 3565 10920 3575
rect 10890 3485 10895 3565
rect 10915 3485 10920 3565
rect 10890 3475 10920 3485
rect 10980 3565 11010 3575
rect 10980 3485 10985 3565
rect 11005 3485 11010 3565
rect 10980 3475 11010 3485
rect 11070 3565 11100 3575
rect 11070 3485 11075 3565
rect 11095 3485 11100 3565
rect 11070 3475 11100 3485
rect 11160 3565 11190 3575
rect 11160 3485 11165 3565
rect 11185 3485 11190 3565
rect 11160 3475 11190 3485
rect 11250 3565 11280 3575
rect 11250 3485 11255 3565
rect 11275 3485 11280 3565
rect 11250 3475 11280 3485
rect 11340 3565 11370 3575
rect 11340 3485 11345 3565
rect 11365 3485 11370 3565
rect 11340 3475 11370 3485
rect 11430 3565 11460 3575
rect 11430 3485 11435 3565
rect 11455 3485 11460 3565
rect 11430 3475 11460 3485
rect 11520 3565 11550 3575
rect 11520 3485 11525 3565
rect 11545 3485 11550 3565
rect 11520 3475 11550 3485
rect 11610 3565 11640 3575
rect 11610 3485 11615 3565
rect 11635 3485 11640 3565
rect 11610 3475 11640 3485
rect 11700 3565 11730 3575
rect 11700 3485 11705 3565
rect 11725 3485 11730 3565
rect 11700 3475 11730 3485
rect 11790 3565 11820 3575
rect 11790 3485 11795 3565
rect 11815 3485 11820 3565
rect 11790 3475 11820 3485
rect 11880 3565 11910 3575
rect 11880 3485 11885 3565
rect 11905 3485 11910 3565
rect 11880 3475 11910 3485
rect 11970 3565 12000 3575
rect 11970 3485 11975 3565
rect 11995 3485 12000 3565
rect 11970 3475 12000 3485
rect 12060 3565 12090 3575
rect 12060 3485 12065 3565
rect 12085 3485 12090 3565
rect 12060 3475 12090 3485
rect 12150 3565 12180 3575
rect 12150 3485 12155 3565
rect 12175 3485 12180 3565
rect 12150 3475 12180 3485
rect 12240 3565 12270 3575
rect 12240 3485 12245 3565
rect 12265 3485 12270 3565
rect 12240 3475 12270 3485
rect 12330 3565 12360 3575
rect 12330 3485 12335 3565
rect 12355 3485 12360 3565
rect 12330 3475 12360 3485
rect 12420 3565 12450 3575
rect 12420 3485 12425 3565
rect 12445 3485 12450 3565
rect 12420 3475 12450 3485
rect 12510 3565 12540 3575
rect 12510 3485 12515 3565
rect 12535 3485 12540 3565
rect 12510 3475 12540 3485
rect 12600 3565 12630 3575
rect 12600 3485 12605 3565
rect 12625 3485 12630 3565
rect 12600 3475 12630 3485
rect 12690 3565 12720 3575
rect 12690 3485 12695 3565
rect 12715 3485 12720 3565
rect 12690 3475 12720 3485
rect 12780 3565 12810 3575
rect 12780 3485 12785 3565
rect 12805 3485 12810 3565
rect 12780 3475 12810 3485
rect 12870 3565 12900 3575
rect 12870 3485 12875 3565
rect 12895 3485 12900 3565
rect 12870 3475 12900 3485
rect 12960 3565 12990 3575
rect 12960 3485 12965 3565
rect 12985 3485 12990 3565
rect 12960 3475 12990 3485
rect 13050 3565 13080 3575
rect 13050 3485 13055 3565
rect 13075 3485 13080 3565
rect 13050 3475 13080 3485
rect 13140 3565 13170 3575
rect 13140 3485 13145 3565
rect 13165 3485 13170 3565
rect 13140 3475 13170 3485
rect 13230 3565 13260 3575
rect 13230 3485 13235 3565
rect 13255 3485 13260 3565
rect 13230 3475 13260 3485
rect 13320 3565 13350 3575
rect 13320 3485 13325 3565
rect 13345 3485 13350 3565
rect 13320 3475 13350 3485
rect 13410 3565 13440 3575
rect 13410 3485 13415 3565
rect 13435 3485 13440 3565
rect 13410 3475 13440 3485
rect 13500 3565 13530 3575
rect 13500 3485 13505 3565
rect 13525 3485 13530 3565
rect 13500 3475 13530 3485
rect 13590 3565 13620 3575
rect 13590 3485 13595 3565
rect 13615 3485 13620 3565
rect 13590 3475 13620 3485
rect 13680 3565 13710 3575
rect 13680 3485 13685 3565
rect 13705 3485 13710 3565
rect 13680 3475 13710 3485
rect 13770 3565 13800 3575
rect 13770 3485 13775 3565
rect 13795 3485 13800 3565
rect 13770 3475 13800 3485
rect 13860 3565 13890 3575
rect 13860 3485 13865 3565
rect 13885 3485 13890 3565
rect 13860 3475 13890 3485
rect 13950 3565 13980 3575
rect 13950 3485 13955 3565
rect 13975 3485 13980 3565
rect 13950 3475 13980 3485
rect 14040 3565 14070 3575
rect 14040 3485 14045 3565
rect 14065 3485 14070 3565
rect 14040 3475 14070 3485
rect 14130 3565 14160 3575
rect 14130 3485 14135 3565
rect 14155 3485 14160 3565
rect 14130 3475 14160 3485
rect 14220 3565 14250 3575
rect 14220 3485 14225 3565
rect 14245 3485 14250 3565
rect 14220 3475 14250 3485
rect 14310 3565 14340 3575
rect 14310 3485 14315 3565
rect 14335 3485 14340 3565
rect 14310 3475 14340 3485
rect 14400 3565 14430 3575
rect 14400 3485 14405 3565
rect 14425 3485 14430 3565
rect 14400 3475 14430 3485
rect 14490 3565 14520 3575
rect 14490 3485 14495 3565
rect 14515 3485 14520 3565
rect 14490 3475 14520 3485
rect 14580 3565 14610 3575
rect 14580 3485 14585 3565
rect 14605 3485 14610 3565
rect 14580 3475 14610 3485
rect 14670 3565 14700 3575
rect 14670 3485 14675 3565
rect 14695 3485 14700 3565
rect 14670 3475 14700 3485
rect 14760 3565 14790 3575
rect 14760 3485 14765 3565
rect 14785 3485 14790 3565
rect 14760 3475 14790 3485
rect 14850 3565 14880 3575
rect 14850 3485 14855 3565
rect 14875 3485 14880 3565
rect 14850 3475 14880 3485
rect 14940 3565 14970 3575
rect 14940 3485 14945 3565
rect 14965 3485 14970 3565
rect 14940 3475 14970 3485
rect 15030 3565 15060 3575
rect 15030 3485 15035 3565
rect 15055 3485 15060 3565
rect 15030 3475 15060 3485
rect 15120 3565 15150 3575
rect 15120 3485 15125 3565
rect 15145 3485 15150 3565
rect 15120 3475 15150 3485
rect 15210 3565 15240 3575
rect 15210 3485 15215 3565
rect 15235 3485 15240 3565
rect 15210 3475 15240 3485
rect 15300 3565 15330 3575
rect 15300 3485 15305 3565
rect 15325 3485 15330 3565
rect 15300 3475 15330 3485
rect 15390 3565 15420 3575
rect 15390 3485 15395 3565
rect 15415 3485 15420 3565
rect 15390 3475 15420 3485
rect 15480 3565 15510 3575
rect 15480 3485 15485 3565
rect 15505 3485 15510 3565
rect 15480 3475 15510 3485
rect 15570 3565 15600 3575
rect 15570 3485 15575 3565
rect 15595 3485 15600 3565
rect 15570 3475 15600 3485
rect 15660 3565 15690 3575
rect 15660 3485 15665 3565
rect 15685 3485 15690 3565
rect 15660 3475 15690 3485
rect 15750 3565 15780 3575
rect 15750 3485 15755 3565
rect 15775 3485 15780 3565
rect 15750 3475 15780 3485
rect 15840 3565 15870 3575
rect 15840 3485 15845 3565
rect 15865 3485 15870 3565
rect 15840 3475 15870 3485
rect 15930 3565 15960 3575
rect 15930 3485 15935 3565
rect 15955 3485 15960 3565
rect 15930 3475 15960 3485
rect 16020 3565 16050 3575
rect 16020 3485 16025 3565
rect 16045 3485 16050 3565
rect 16020 3475 16050 3485
rect 16110 3565 16140 3575
rect 16110 3485 16115 3565
rect 16135 3485 16140 3565
rect 16110 3475 16140 3485
rect 16200 3565 16230 3575
rect 16200 3485 16205 3565
rect 16225 3485 16230 3565
rect 16200 3475 16230 3485
rect 16290 3565 16320 3575
rect 16290 3485 16295 3565
rect 16315 3485 16320 3565
rect 16290 3475 16320 3485
rect 16380 3565 16410 3575
rect 16380 3485 16385 3565
rect 16405 3485 16410 3565
rect 16380 3475 16410 3485
rect 16470 3565 16500 3575
rect 16470 3485 16475 3565
rect 16495 3485 16500 3565
rect 16470 3475 16500 3485
rect 16560 3565 16590 3575
rect 16560 3485 16565 3565
rect 16585 3485 16590 3565
rect 16560 3475 16590 3485
rect 16650 3565 16680 3575
rect 16650 3485 16655 3565
rect 16675 3485 16680 3565
rect 16650 3475 16680 3485
rect 16740 3565 16770 3575
rect 16740 3485 16745 3565
rect 16765 3485 16770 3565
rect 16740 3475 16770 3485
rect 16830 3565 16860 3575
rect 16830 3485 16835 3565
rect 16855 3485 16860 3565
rect 16830 3475 16860 3485
rect 16920 3565 16950 3575
rect 16920 3485 16925 3565
rect 16945 3485 16950 3565
rect 16920 3475 16950 3485
rect 17010 3565 17040 3575
rect 17010 3485 17015 3565
rect 17035 3485 17040 3565
rect 17010 3475 17040 3485
rect 17100 3565 17130 3575
rect 17100 3485 17105 3565
rect 17125 3485 17130 3565
rect 17100 3475 17130 3485
rect 17190 3565 17220 3575
rect 17190 3485 17195 3565
rect 17215 3485 17220 3565
rect 17190 3475 17220 3485
rect 17280 3565 17310 3575
rect 17280 3485 17285 3565
rect 17305 3485 17310 3565
rect 17280 3475 17310 3485
rect 17370 3565 17400 3575
rect 17370 3485 17375 3565
rect 17395 3485 17400 3565
rect 17370 3475 17400 3485
rect 17460 3565 17490 3575
rect 17460 3485 17465 3565
rect 17485 3485 17490 3565
rect 17460 3475 17490 3485
rect 17550 3565 17580 3575
rect 17550 3485 17555 3565
rect 17575 3485 17580 3565
rect 17550 3475 17580 3485
rect 17640 3565 17670 3575
rect 17640 3485 17645 3565
rect 17665 3485 17670 3565
rect 17640 3475 17670 3485
rect 17730 3565 17760 3575
rect 17730 3485 17735 3565
rect 17755 3485 17760 3565
rect 17730 3475 17760 3485
rect 17820 3565 17850 3575
rect 17820 3485 17825 3565
rect 17845 3485 17850 3565
rect 17820 3475 17850 3485
rect 17910 3565 17940 3575
rect 17910 3485 17915 3565
rect 17935 3485 17940 3565
rect 17910 3475 17940 3485
rect 18000 3565 18030 3575
rect 18000 3485 18005 3565
rect 18025 3485 18030 3565
rect 18000 3475 18030 3485
rect 18090 3565 18120 3575
rect 18090 3485 18095 3565
rect 18115 3485 18120 3565
rect 18090 3475 18120 3485
rect 18180 3565 18210 3575
rect 18180 3485 18185 3565
rect 18205 3485 18210 3565
rect 18180 3475 18210 3485
rect 18270 3565 18300 3575
rect 18270 3485 18275 3565
rect 18295 3485 18300 3565
rect 18270 3475 18300 3485
rect 18360 3565 18390 3575
rect 18360 3485 18365 3565
rect 18385 3485 18390 3565
rect 18360 3475 18390 3485
rect 18450 3565 18480 3575
rect 18450 3485 18455 3565
rect 18475 3485 18480 3565
rect 18450 3475 18480 3485
rect 18540 3565 18570 3575
rect 18540 3485 18545 3565
rect 18565 3485 18570 3565
rect 18540 3475 18570 3485
rect 18630 3565 18660 3575
rect 18630 3485 18635 3565
rect 18655 3485 18660 3565
rect 18630 3475 18660 3485
rect 18720 3565 18750 3575
rect 18720 3485 18725 3565
rect 18745 3485 18750 3565
rect 18720 3475 18750 3485
rect 18810 3565 18840 3575
rect 18810 3485 18815 3565
rect 18835 3485 18840 3565
rect 18810 3475 18840 3485
rect 18900 3565 18930 3575
rect 18900 3485 18905 3565
rect 18925 3485 18930 3565
rect 18900 3475 18930 3485
rect 18990 3565 19020 3575
rect 18990 3485 18995 3565
rect 19015 3485 19020 3565
rect 18990 3475 19020 3485
rect 19080 3565 19110 3575
rect 19080 3485 19085 3565
rect 19105 3485 19110 3565
rect 19080 3475 19110 3485
rect 19170 3565 19200 3575
rect 19170 3485 19175 3565
rect 19195 3485 19200 3565
rect 19170 3475 19200 3485
rect 19260 3565 19290 3575
rect 19260 3485 19265 3565
rect 19285 3485 19290 3565
rect 19260 3475 19290 3485
rect 19350 3565 19380 3575
rect 19350 3485 19355 3565
rect 19375 3485 19380 3565
rect 19350 3475 19380 3485
rect 19440 3565 19470 3575
rect 19440 3485 19445 3565
rect 19465 3485 19470 3565
rect 19440 3475 19470 3485
rect 19530 3565 19560 3575
rect 19530 3485 19535 3565
rect 19555 3485 19560 3565
rect 19530 3475 19560 3485
rect 19620 3565 19650 3575
rect 19620 3485 19625 3565
rect 19645 3485 19650 3565
rect 19620 3475 19650 3485
rect 19710 3565 19740 3575
rect 19710 3485 19715 3565
rect 19735 3485 19740 3565
rect 19710 3475 19740 3485
rect 19800 3565 19830 3575
rect 19800 3485 19805 3565
rect 19825 3485 19830 3565
rect 19800 3475 19830 3485
rect 19890 3565 19920 3575
rect 19890 3485 19895 3565
rect 19915 3485 19920 3565
rect 19890 3475 19920 3485
rect 19980 3565 20010 3575
rect 19980 3485 19985 3565
rect 20005 3485 20010 3565
rect 19980 3475 20010 3485
rect 20070 3475 20100 3575
rect 20160 3475 20190 3575
rect 20250 3475 20280 3575
rect 20340 3475 20370 3575
rect 20430 3475 20460 3575
rect 20520 3475 20550 3575
rect 20610 3475 20640 3575
rect 20700 3565 20730 3575
rect 20700 3485 20705 3565
rect 20725 3485 20730 3565
rect 20700 3475 20730 3485
rect 9185 3455 9205 3475
rect 9905 3455 9925 3475
rect 10625 3455 10645 3475
rect 11345 3455 11365 3475
rect 12065 3455 12085 3475
rect 12785 3455 12805 3475
rect 13505 3455 13525 3475
rect 14225 3455 14245 3475
rect 14945 3455 14965 3475
rect 15665 3455 15685 3475
rect 16385 3455 16405 3475
rect 17105 3455 17125 3475
rect 17825 3455 17845 3475
rect 18545 3455 18565 3475
rect 19265 3455 19285 3475
rect 19985 3455 20005 3475
rect 20705 3455 20725 3475
rect 9040 3420 9045 3450
rect 9075 3420 9080 3450
rect 9040 3415 9080 3420
rect 9175 3450 9215 3455
rect 9175 3420 9180 3450
rect 9210 3420 9215 3450
rect 9175 3415 9215 3420
rect 9895 3450 9935 3455
rect 9895 3420 9900 3450
rect 9930 3420 9935 3450
rect 9895 3415 9935 3420
rect 10075 3450 10115 3455
rect 10075 3420 10080 3450
rect 10110 3420 10115 3450
rect 10075 3415 10115 3420
rect 10255 3450 10295 3455
rect 10255 3420 10260 3450
rect 10290 3420 10295 3450
rect 10255 3415 10295 3420
rect 10435 3450 10475 3455
rect 10435 3420 10440 3450
rect 10470 3420 10475 3450
rect 10435 3415 10475 3420
rect 10615 3450 10655 3455
rect 10615 3420 10620 3450
rect 10650 3420 10655 3450
rect 10615 3415 10655 3420
rect 10795 3450 10835 3455
rect 10795 3420 10800 3450
rect 10830 3420 10835 3450
rect 10795 3415 10835 3420
rect 10975 3450 11015 3455
rect 10975 3420 10980 3450
rect 11010 3420 11015 3450
rect 10975 3415 11015 3420
rect 11155 3450 11195 3455
rect 11155 3420 11160 3450
rect 11190 3420 11195 3450
rect 11155 3415 11195 3420
rect 11335 3450 11375 3455
rect 11335 3420 11340 3450
rect 11370 3420 11375 3450
rect 11335 3415 11375 3420
rect 11515 3450 11555 3455
rect 11515 3420 11520 3450
rect 11550 3420 11555 3450
rect 11515 3415 11555 3420
rect 11695 3450 11735 3455
rect 11695 3420 11700 3450
rect 11730 3420 11735 3450
rect 11695 3415 11735 3420
rect 11875 3450 11915 3455
rect 11875 3420 11880 3450
rect 11910 3420 11915 3450
rect 11875 3415 11915 3420
rect 12055 3450 12095 3455
rect 12055 3420 12060 3450
rect 12090 3420 12095 3450
rect 12055 3415 12095 3420
rect 12235 3450 12275 3455
rect 12235 3420 12240 3450
rect 12270 3420 12275 3450
rect 12235 3415 12275 3420
rect 12415 3450 12455 3455
rect 12415 3420 12420 3450
rect 12450 3420 12455 3450
rect 12415 3415 12455 3420
rect 12595 3450 12635 3455
rect 12595 3420 12600 3450
rect 12630 3420 12635 3450
rect 12595 3415 12635 3420
rect 12775 3450 12815 3455
rect 12775 3420 12780 3450
rect 12810 3420 12815 3450
rect 12775 3415 12815 3420
rect 12955 3450 12995 3455
rect 12955 3420 12960 3450
rect 12990 3420 12995 3450
rect 12955 3415 12995 3420
rect 13135 3450 13175 3455
rect 13135 3420 13140 3450
rect 13170 3420 13175 3450
rect 13135 3415 13175 3420
rect 13315 3450 13355 3455
rect 13315 3420 13320 3450
rect 13350 3420 13355 3450
rect 13315 3415 13355 3420
rect 13495 3450 13535 3455
rect 13495 3420 13500 3450
rect 13530 3420 13535 3450
rect 13495 3415 13535 3420
rect 13675 3450 13715 3455
rect 13675 3420 13680 3450
rect 13710 3420 13715 3450
rect 13675 3415 13715 3420
rect 13855 3450 13895 3455
rect 13855 3420 13860 3450
rect 13890 3420 13895 3450
rect 13855 3415 13895 3420
rect 14035 3450 14075 3455
rect 14035 3420 14040 3450
rect 14070 3420 14075 3450
rect 14035 3415 14075 3420
rect 14215 3450 14255 3455
rect 14215 3420 14220 3450
rect 14250 3420 14255 3450
rect 14215 3415 14255 3420
rect 14395 3450 14435 3455
rect 14395 3420 14400 3450
rect 14430 3420 14435 3450
rect 14395 3415 14435 3420
rect 14575 3450 14615 3455
rect 14575 3420 14580 3450
rect 14610 3420 14615 3450
rect 14575 3415 14615 3420
rect 14755 3450 14795 3455
rect 14755 3420 14760 3450
rect 14790 3420 14795 3450
rect 14755 3415 14795 3420
rect 14935 3450 14975 3455
rect 14935 3420 14940 3450
rect 14970 3420 14975 3450
rect 14935 3415 14975 3420
rect 15115 3450 15155 3455
rect 15115 3420 15120 3450
rect 15150 3420 15155 3450
rect 15115 3415 15155 3420
rect 15295 3450 15335 3455
rect 15295 3420 15300 3450
rect 15330 3420 15335 3450
rect 15295 3415 15335 3420
rect 15475 3450 15515 3455
rect 15475 3420 15480 3450
rect 15510 3420 15515 3450
rect 15475 3415 15515 3420
rect 15655 3450 15695 3455
rect 15655 3420 15660 3450
rect 15690 3420 15695 3450
rect 15655 3415 15695 3420
rect 15835 3450 15875 3455
rect 15835 3420 15840 3450
rect 15870 3420 15875 3450
rect 15835 3415 15875 3420
rect 16015 3450 16055 3455
rect 16015 3420 16020 3450
rect 16050 3420 16055 3450
rect 16015 3415 16055 3420
rect 16195 3450 16235 3455
rect 16195 3420 16200 3450
rect 16230 3420 16235 3450
rect 16195 3415 16235 3420
rect 16375 3450 16415 3455
rect 16375 3420 16380 3450
rect 16410 3420 16415 3450
rect 16375 3415 16415 3420
rect 16555 3450 16595 3455
rect 16555 3420 16560 3450
rect 16590 3420 16595 3450
rect 16555 3415 16595 3420
rect 16735 3450 16775 3455
rect 16735 3420 16740 3450
rect 16770 3420 16775 3450
rect 16735 3415 16775 3420
rect 16915 3450 16955 3455
rect 16915 3420 16920 3450
rect 16950 3420 16955 3450
rect 16915 3415 16955 3420
rect 17095 3450 17135 3455
rect 17095 3420 17100 3450
rect 17130 3420 17135 3450
rect 17095 3415 17135 3420
rect 17275 3450 17315 3455
rect 17275 3420 17280 3450
rect 17310 3420 17315 3450
rect 17275 3415 17315 3420
rect 17455 3450 17495 3455
rect 17455 3420 17460 3450
rect 17490 3420 17495 3450
rect 17455 3415 17495 3420
rect 17635 3450 17675 3455
rect 17635 3420 17640 3450
rect 17670 3420 17675 3450
rect 17635 3415 17675 3420
rect 17815 3450 17855 3455
rect 17815 3420 17820 3450
rect 17850 3420 17855 3450
rect 17815 3415 17855 3420
rect 17995 3450 18035 3455
rect 17995 3420 18000 3450
rect 18030 3420 18035 3450
rect 17995 3415 18035 3420
rect 18175 3450 18215 3455
rect 18175 3420 18180 3450
rect 18210 3420 18215 3450
rect 18175 3415 18215 3420
rect 18355 3450 18395 3455
rect 18355 3420 18360 3450
rect 18390 3420 18395 3450
rect 18355 3415 18395 3420
rect 18535 3450 18575 3455
rect 18535 3420 18540 3450
rect 18570 3420 18575 3450
rect 18535 3415 18575 3420
rect 18715 3450 18755 3455
rect 18715 3420 18720 3450
rect 18750 3420 18755 3450
rect 18715 3415 18755 3420
rect 18895 3450 18935 3455
rect 18895 3420 18900 3450
rect 18930 3420 18935 3450
rect 18895 3415 18935 3420
rect 19075 3450 19115 3455
rect 19075 3420 19080 3450
rect 19110 3420 19115 3450
rect 19075 3415 19115 3420
rect 19255 3450 19295 3455
rect 19255 3420 19260 3450
rect 19290 3420 19295 3450
rect 19255 3415 19295 3420
rect 19435 3450 19475 3455
rect 19435 3420 19440 3450
rect 19470 3420 19475 3450
rect 19435 3415 19475 3420
rect 19615 3450 19655 3455
rect 19615 3420 19620 3450
rect 19650 3420 19655 3450
rect 19615 3415 19655 3420
rect 19795 3450 19835 3455
rect 19795 3420 19800 3450
rect 19830 3420 19835 3450
rect 19795 3415 19835 3420
rect 19975 3450 20015 3455
rect 19975 3420 19980 3450
rect 20010 3420 20015 3450
rect 19975 3415 20015 3420
rect 20695 3450 20735 3455
rect 20695 3420 20700 3450
rect 20730 3420 20735 3450
rect 20695 3415 20735 3420
rect 20830 3450 20870 4375
rect 20830 3420 20835 3450
rect 20865 3420 20870 3450
rect 20830 3415 20870 3420
<< via1 >>
rect 9180 4365 9210 4370
rect 9180 4345 9185 4365
rect 9185 4345 9205 4365
rect 9205 4345 9210 4365
rect 9180 4340 9210 4345
rect 9900 4365 9930 4370
rect 9900 4345 9905 4365
rect 9905 4345 9925 4365
rect 9925 4345 9930 4365
rect 9900 4340 9930 4345
rect 10080 4365 10110 4370
rect 10080 4345 10085 4365
rect 10085 4345 10105 4365
rect 10105 4345 10110 4365
rect 10080 4340 10110 4345
rect 10260 4365 10290 4370
rect 10260 4345 10265 4365
rect 10265 4345 10285 4365
rect 10285 4345 10290 4365
rect 10260 4340 10290 4345
rect 10440 4365 10470 4370
rect 10440 4345 10445 4365
rect 10445 4345 10465 4365
rect 10465 4345 10470 4365
rect 10440 4340 10470 4345
rect 10620 4365 10650 4370
rect 10620 4345 10625 4365
rect 10625 4345 10645 4365
rect 10645 4345 10650 4365
rect 10620 4340 10650 4345
rect 10800 4365 10830 4370
rect 10800 4345 10805 4365
rect 10805 4345 10825 4365
rect 10825 4345 10830 4365
rect 10800 4340 10830 4345
rect 10980 4365 11010 4370
rect 10980 4345 10985 4365
rect 10985 4345 11005 4365
rect 11005 4345 11010 4365
rect 10980 4340 11010 4345
rect 11160 4365 11190 4370
rect 11160 4345 11165 4365
rect 11165 4345 11185 4365
rect 11185 4345 11190 4365
rect 11160 4340 11190 4345
rect 11340 4365 11370 4370
rect 11340 4345 11345 4365
rect 11345 4345 11365 4365
rect 11365 4345 11370 4365
rect 11340 4340 11370 4345
rect 11520 4365 11550 4370
rect 11520 4345 11525 4365
rect 11525 4345 11545 4365
rect 11545 4345 11550 4365
rect 11520 4340 11550 4345
rect 11700 4365 11730 4370
rect 11700 4345 11705 4365
rect 11705 4345 11725 4365
rect 11725 4345 11730 4365
rect 11700 4340 11730 4345
rect 11880 4365 11910 4370
rect 11880 4345 11885 4365
rect 11885 4345 11905 4365
rect 11905 4345 11910 4365
rect 11880 4340 11910 4345
rect 12060 4365 12090 4370
rect 12060 4345 12065 4365
rect 12065 4345 12085 4365
rect 12085 4345 12090 4365
rect 12060 4340 12090 4345
rect 12240 4365 12270 4370
rect 12240 4345 12245 4365
rect 12245 4345 12265 4365
rect 12265 4345 12270 4365
rect 12240 4340 12270 4345
rect 12420 4365 12450 4370
rect 12420 4345 12425 4365
rect 12425 4345 12445 4365
rect 12445 4345 12450 4365
rect 12420 4340 12450 4345
rect 12600 4365 12630 4370
rect 12600 4345 12605 4365
rect 12605 4345 12625 4365
rect 12625 4345 12630 4365
rect 12600 4340 12630 4345
rect 12780 4365 12810 4370
rect 12780 4345 12785 4365
rect 12785 4345 12805 4365
rect 12805 4345 12810 4365
rect 12780 4340 12810 4345
rect 12960 4365 12990 4370
rect 12960 4345 12965 4365
rect 12965 4345 12985 4365
rect 12985 4345 12990 4365
rect 12960 4340 12990 4345
rect 13140 4365 13170 4370
rect 13140 4345 13145 4365
rect 13145 4345 13165 4365
rect 13165 4345 13170 4365
rect 13140 4340 13170 4345
rect 13320 4365 13350 4370
rect 13320 4345 13325 4365
rect 13325 4345 13345 4365
rect 13345 4345 13350 4365
rect 13320 4340 13350 4345
rect 13500 4365 13530 4370
rect 13500 4345 13505 4365
rect 13505 4345 13525 4365
rect 13525 4345 13530 4365
rect 13500 4340 13530 4345
rect 13680 4365 13710 4370
rect 13680 4345 13685 4365
rect 13685 4345 13705 4365
rect 13705 4345 13710 4365
rect 13680 4340 13710 4345
rect 13860 4365 13890 4370
rect 13860 4345 13865 4365
rect 13865 4345 13885 4365
rect 13885 4345 13890 4365
rect 13860 4340 13890 4345
rect 14040 4365 14070 4370
rect 14040 4345 14045 4365
rect 14045 4345 14065 4365
rect 14065 4345 14070 4365
rect 14040 4340 14070 4345
rect 14220 4365 14250 4370
rect 14220 4345 14225 4365
rect 14225 4345 14245 4365
rect 14245 4345 14250 4365
rect 14220 4340 14250 4345
rect 14400 4365 14430 4370
rect 14400 4345 14405 4365
rect 14405 4345 14425 4365
rect 14425 4345 14430 4365
rect 14400 4340 14430 4345
rect 14580 4365 14610 4370
rect 14580 4345 14585 4365
rect 14585 4345 14605 4365
rect 14605 4345 14610 4365
rect 14580 4340 14610 4345
rect 14760 4365 14790 4370
rect 14760 4345 14765 4365
rect 14765 4345 14785 4365
rect 14785 4345 14790 4365
rect 14760 4340 14790 4345
rect 14940 4365 14970 4370
rect 14940 4345 14945 4365
rect 14945 4345 14965 4365
rect 14965 4345 14970 4365
rect 14940 4340 14970 4345
rect 15120 4365 15150 4370
rect 15120 4345 15125 4365
rect 15125 4345 15145 4365
rect 15145 4345 15150 4365
rect 15120 4340 15150 4345
rect 15300 4365 15330 4370
rect 15300 4345 15305 4365
rect 15305 4345 15325 4365
rect 15325 4345 15330 4365
rect 15300 4340 15330 4345
rect 15480 4365 15510 4370
rect 15480 4345 15485 4365
rect 15485 4345 15505 4365
rect 15505 4345 15510 4365
rect 15480 4340 15510 4345
rect 15660 4365 15690 4370
rect 15660 4345 15665 4365
rect 15665 4345 15685 4365
rect 15685 4345 15690 4365
rect 15660 4340 15690 4345
rect 15840 4365 15870 4370
rect 15840 4345 15845 4365
rect 15845 4345 15865 4365
rect 15865 4345 15870 4365
rect 15840 4340 15870 4345
rect 16020 4365 16050 4370
rect 16020 4345 16025 4365
rect 16025 4345 16045 4365
rect 16045 4345 16050 4365
rect 16020 4340 16050 4345
rect 16200 4365 16230 4370
rect 16200 4345 16205 4365
rect 16205 4345 16225 4365
rect 16225 4345 16230 4365
rect 16200 4340 16230 4345
rect 16380 4365 16410 4370
rect 16380 4345 16385 4365
rect 16385 4345 16405 4365
rect 16405 4345 16410 4365
rect 16380 4340 16410 4345
rect 16560 4365 16590 4370
rect 16560 4345 16565 4365
rect 16565 4345 16585 4365
rect 16585 4345 16590 4365
rect 16560 4340 16590 4345
rect 16740 4365 16770 4370
rect 16740 4345 16745 4365
rect 16745 4345 16765 4365
rect 16765 4345 16770 4365
rect 16740 4340 16770 4345
rect 16920 4365 16950 4370
rect 16920 4345 16925 4365
rect 16925 4345 16945 4365
rect 16945 4345 16950 4365
rect 16920 4340 16950 4345
rect 17100 4365 17130 4370
rect 17100 4345 17105 4365
rect 17105 4345 17125 4365
rect 17125 4345 17130 4365
rect 17100 4340 17130 4345
rect 17280 4365 17310 4370
rect 17280 4345 17285 4365
rect 17285 4345 17305 4365
rect 17305 4345 17310 4365
rect 17280 4340 17310 4345
rect 17460 4365 17490 4370
rect 17460 4345 17465 4365
rect 17465 4345 17485 4365
rect 17485 4345 17490 4365
rect 17460 4340 17490 4345
rect 17640 4365 17670 4370
rect 17640 4345 17645 4365
rect 17645 4345 17665 4365
rect 17665 4345 17670 4365
rect 17640 4340 17670 4345
rect 17820 4365 17850 4370
rect 17820 4345 17825 4365
rect 17825 4345 17845 4365
rect 17845 4345 17850 4365
rect 17820 4340 17850 4345
rect 18000 4365 18030 4370
rect 18000 4345 18005 4365
rect 18005 4345 18025 4365
rect 18025 4345 18030 4365
rect 18000 4340 18030 4345
rect 18180 4365 18210 4370
rect 18180 4345 18185 4365
rect 18185 4345 18205 4365
rect 18205 4345 18210 4365
rect 18180 4340 18210 4345
rect 18360 4365 18390 4370
rect 18360 4345 18365 4365
rect 18365 4345 18385 4365
rect 18385 4345 18390 4365
rect 18360 4340 18390 4345
rect 18540 4365 18570 4370
rect 18540 4345 18545 4365
rect 18545 4345 18565 4365
rect 18565 4345 18570 4365
rect 18540 4340 18570 4345
rect 18720 4365 18750 4370
rect 18720 4345 18725 4365
rect 18725 4345 18745 4365
rect 18745 4345 18750 4365
rect 18720 4340 18750 4345
rect 18900 4365 18930 4370
rect 18900 4345 18905 4365
rect 18905 4345 18925 4365
rect 18925 4345 18930 4365
rect 18900 4340 18930 4345
rect 19080 4365 19110 4370
rect 19080 4345 19085 4365
rect 19085 4345 19105 4365
rect 19105 4345 19110 4365
rect 19080 4340 19110 4345
rect 19260 4365 19290 4370
rect 19260 4345 19265 4365
rect 19265 4345 19285 4365
rect 19285 4345 19290 4365
rect 19260 4340 19290 4345
rect 19440 4365 19470 4370
rect 19440 4345 19445 4365
rect 19445 4345 19465 4365
rect 19465 4345 19470 4365
rect 19440 4340 19470 4345
rect 19620 4365 19650 4370
rect 19620 4345 19625 4365
rect 19625 4345 19645 4365
rect 19645 4345 19650 4365
rect 19620 4340 19650 4345
rect 19800 4365 19830 4370
rect 19800 4345 19805 4365
rect 19805 4345 19825 4365
rect 19825 4345 19830 4365
rect 19800 4340 19830 4345
rect 19980 4365 20010 4370
rect 19980 4345 19985 4365
rect 19985 4345 20005 4365
rect 20005 4345 20010 4365
rect 19980 4340 20010 4345
rect 20700 4365 20730 4370
rect 20700 4345 20705 4365
rect 20705 4345 20725 4365
rect 20725 4345 20730 4365
rect 20700 4340 20730 4345
rect 9045 3445 9075 3450
rect 9045 3425 9050 3445
rect 9050 3425 9070 3445
rect 9070 3425 9075 3445
rect 9045 3420 9075 3425
rect 9180 3445 9210 3450
rect 9180 3425 9185 3445
rect 9185 3425 9205 3445
rect 9205 3425 9210 3445
rect 9180 3420 9210 3425
rect 9900 3445 9930 3450
rect 9900 3425 9905 3445
rect 9905 3425 9925 3445
rect 9925 3425 9930 3445
rect 9900 3420 9930 3425
rect 10080 3445 10110 3450
rect 10080 3425 10085 3445
rect 10085 3425 10105 3445
rect 10105 3425 10110 3445
rect 10080 3420 10110 3425
rect 10260 3445 10290 3450
rect 10260 3425 10265 3445
rect 10265 3425 10285 3445
rect 10285 3425 10290 3445
rect 10260 3420 10290 3425
rect 10440 3445 10470 3450
rect 10440 3425 10445 3445
rect 10445 3425 10465 3445
rect 10465 3425 10470 3445
rect 10440 3420 10470 3425
rect 10620 3445 10650 3450
rect 10620 3425 10625 3445
rect 10625 3425 10645 3445
rect 10645 3425 10650 3445
rect 10620 3420 10650 3425
rect 10800 3445 10830 3450
rect 10800 3425 10805 3445
rect 10805 3425 10825 3445
rect 10825 3425 10830 3445
rect 10800 3420 10830 3425
rect 10980 3445 11010 3450
rect 10980 3425 10985 3445
rect 10985 3425 11005 3445
rect 11005 3425 11010 3445
rect 10980 3420 11010 3425
rect 11160 3445 11190 3450
rect 11160 3425 11165 3445
rect 11165 3425 11185 3445
rect 11185 3425 11190 3445
rect 11160 3420 11190 3425
rect 11340 3445 11370 3450
rect 11340 3425 11345 3445
rect 11345 3425 11365 3445
rect 11365 3425 11370 3445
rect 11340 3420 11370 3425
rect 11520 3445 11550 3450
rect 11520 3425 11525 3445
rect 11525 3425 11545 3445
rect 11545 3425 11550 3445
rect 11520 3420 11550 3425
rect 11700 3445 11730 3450
rect 11700 3425 11705 3445
rect 11705 3425 11725 3445
rect 11725 3425 11730 3445
rect 11700 3420 11730 3425
rect 11880 3445 11910 3450
rect 11880 3425 11885 3445
rect 11885 3425 11905 3445
rect 11905 3425 11910 3445
rect 11880 3420 11910 3425
rect 12060 3445 12090 3450
rect 12060 3425 12065 3445
rect 12065 3425 12085 3445
rect 12085 3425 12090 3445
rect 12060 3420 12090 3425
rect 12240 3445 12270 3450
rect 12240 3425 12245 3445
rect 12245 3425 12265 3445
rect 12265 3425 12270 3445
rect 12240 3420 12270 3425
rect 12420 3445 12450 3450
rect 12420 3425 12425 3445
rect 12425 3425 12445 3445
rect 12445 3425 12450 3445
rect 12420 3420 12450 3425
rect 12600 3445 12630 3450
rect 12600 3425 12605 3445
rect 12605 3425 12625 3445
rect 12625 3425 12630 3445
rect 12600 3420 12630 3425
rect 12780 3445 12810 3450
rect 12780 3425 12785 3445
rect 12785 3425 12805 3445
rect 12805 3425 12810 3445
rect 12780 3420 12810 3425
rect 12960 3445 12990 3450
rect 12960 3425 12965 3445
rect 12965 3425 12985 3445
rect 12985 3425 12990 3445
rect 12960 3420 12990 3425
rect 13140 3445 13170 3450
rect 13140 3425 13145 3445
rect 13145 3425 13165 3445
rect 13165 3425 13170 3445
rect 13140 3420 13170 3425
rect 13320 3445 13350 3450
rect 13320 3425 13325 3445
rect 13325 3425 13345 3445
rect 13345 3425 13350 3445
rect 13320 3420 13350 3425
rect 13500 3445 13530 3450
rect 13500 3425 13505 3445
rect 13505 3425 13525 3445
rect 13525 3425 13530 3445
rect 13500 3420 13530 3425
rect 13680 3445 13710 3450
rect 13680 3425 13685 3445
rect 13685 3425 13705 3445
rect 13705 3425 13710 3445
rect 13680 3420 13710 3425
rect 13860 3445 13890 3450
rect 13860 3425 13865 3445
rect 13865 3425 13885 3445
rect 13885 3425 13890 3445
rect 13860 3420 13890 3425
rect 14040 3445 14070 3450
rect 14040 3425 14045 3445
rect 14045 3425 14065 3445
rect 14065 3425 14070 3445
rect 14040 3420 14070 3425
rect 14220 3445 14250 3450
rect 14220 3425 14225 3445
rect 14225 3425 14245 3445
rect 14245 3425 14250 3445
rect 14220 3420 14250 3425
rect 14400 3445 14430 3450
rect 14400 3425 14405 3445
rect 14405 3425 14425 3445
rect 14425 3425 14430 3445
rect 14400 3420 14430 3425
rect 14580 3445 14610 3450
rect 14580 3425 14585 3445
rect 14585 3425 14605 3445
rect 14605 3425 14610 3445
rect 14580 3420 14610 3425
rect 14760 3445 14790 3450
rect 14760 3425 14765 3445
rect 14765 3425 14785 3445
rect 14785 3425 14790 3445
rect 14760 3420 14790 3425
rect 14940 3445 14970 3450
rect 14940 3425 14945 3445
rect 14945 3425 14965 3445
rect 14965 3425 14970 3445
rect 14940 3420 14970 3425
rect 15120 3445 15150 3450
rect 15120 3425 15125 3445
rect 15125 3425 15145 3445
rect 15145 3425 15150 3445
rect 15120 3420 15150 3425
rect 15300 3445 15330 3450
rect 15300 3425 15305 3445
rect 15305 3425 15325 3445
rect 15325 3425 15330 3445
rect 15300 3420 15330 3425
rect 15480 3445 15510 3450
rect 15480 3425 15485 3445
rect 15485 3425 15505 3445
rect 15505 3425 15510 3445
rect 15480 3420 15510 3425
rect 15660 3445 15690 3450
rect 15660 3425 15665 3445
rect 15665 3425 15685 3445
rect 15685 3425 15690 3445
rect 15660 3420 15690 3425
rect 15840 3445 15870 3450
rect 15840 3425 15845 3445
rect 15845 3425 15865 3445
rect 15865 3425 15870 3445
rect 15840 3420 15870 3425
rect 16020 3445 16050 3450
rect 16020 3425 16025 3445
rect 16025 3425 16045 3445
rect 16045 3425 16050 3445
rect 16020 3420 16050 3425
rect 16200 3445 16230 3450
rect 16200 3425 16205 3445
rect 16205 3425 16225 3445
rect 16225 3425 16230 3445
rect 16200 3420 16230 3425
rect 16380 3445 16410 3450
rect 16380 3425 16385 3445
rect 16385 3425 16405 3445
rect 16405 3425 16410 3445
rect 16380 3420 16410 3425
rect 16560 3445 16590 3450
rect 16560 3425 16565 3445
rect 16565 3425 16585 3445
rect 16585 3425 16590 3445
rect 16560 3420 16590 3425
rect 16740 3445 16770 3450
rect 16740 3425 16745 3445
rect 16745 3425 16765 3445
rect 16765 3425 16770 3445
rect 16740 3420 16770 3425
rect 16920 3445 16950 3450
rect 16920 3425 16925 3445
rect 16925 3425 16945 3445
rect 16945 3425 16950 3445
rect 16920 3420 16950 3425
rect 17100 3445 17130 3450
rect 17100 3425 17105 3445
rect 17105 3425 17125 3445
rect 17125 3425 17130 3445
rect 17100 3420 17130 3425
rect 17280 3445 17310 3450
rect 17280 3425 17285 3445
rect 17285 3425 17305 3445
rect 17305 3425 17310 3445
rect 17280 3420 17310 3425
rect 17460 3445 17490 3450
rect 17460 3425 17465 3445
rect 17465 3425 17485 3445
rect 17485 3425 17490 3445
rect 17460 3420 17490 3425
rect 17640 3445 17670 3450
rect 17640 3425 17645 3445
rect 17645 3425 17665 3445
rect 17665 3425 17670 3445
rect 17640 3420 17670 3425
rect 17820 3445 17850 3450
rect 17820 3425 17825 3445
rect 17825 3425 17845 3445
rect 17845 3425 17850 3445
rect 17820 3420 17850 3425
rect 18000 3445 18030 3450
rect 18000 3425 18005 3445
rect 18005 3425 18025 3445
rect 18025 3425 18030 3445
rect 18000 3420 18030 3425
rect 18180 3445 18210 3450
rect 18180 3425 18185 3445
rect 18185 3425 18205 3445
rect 18205 3425 18210 3445
rect 18180 3420 18210 3425
rect 18360 3445 18390 3450
rect 18360 3425 18365 3445
rect 18365 3425 18385 3445
rect 18385 3425 18390 3445
rect 18360 3420 18390 3425
rect 18540 3445 18570 3450
rect 18540 3425 18545 3445
rect 18545 3425 18565 3445
rect 18565 3425 18570 3445
rect 18540 3420 18570 3425
rect 18720 3445 18750 3450
rect 18720 3425 18725 3445
rect 18725 3425 18745 3445
rect 18745 3425 18750 3445
rect 18720 3420 18750 3425
rect 18900 3445 18930 3450
rect 18900 3425 18905 3445
rect 18905 3425 18925 3445
rect 18925 3425 18930 3445
rect 18900 3420 18930 3425
rect 19080 3445 19110 3450
rect 19080 3425 19085 3445
rect 19085 3425 19105 3445
rect 19105 3425 19110 3445
rect 19080 3420 19110 3425
rect 19260 3445 19290 3450
rect 19260 3425 19265 3445
rect 19265 3425 19285 3445
rect 19285 3425 19290 3445
rect 19260 3420 19290 3425
rect 19440 3445 19470 3450
rect 19440 3425 19445 3445
rect 19445 3425 19465 3445
rect 19465 3425 19470 3445
rect 19440 3420 19470 3425
rect 19620 3445 19650 3450
rect 19620 3425 19625 3445
rect 19625 3425 19645 3445
rect 19645 3425 19650 3445
rect 19620 3420 19650 3425
rect 19800 3445 19830 3450
rect 19800 3425 19805 3445
rect 19805 3425 19825 3445
rect 19825 3425 19830 3445
rect 19800 3420 19830 3425
rect 19980 3445 20010 3450
rect 19980 3425 19985 3445
rect 19985 3425 20005 3445
rect 20005 3425 20010 3445
rect 19980 3420 20010 3425
rect 20700 3445 20730 3450
rect 20700 3425 20705 3445
rect 20705 3425 20725 3445
rect 20725 3425 20730 3445
rect 20700 3420 20730 3425
rect 20835 3445 20865 3450
rect 20835 3425 20840 3445
rect 20840 3425 20860 3445
rect 20860 3425 20865 3445
rect 20835 3420 20865 3425
<< metal2 >>
rect 9175 4370 20740 4375
rect 9175 4340 9180 4370
rect 9210 4340 9900 4370
rect 9930 4340 10080 4370
rect 10110 4340 10260 4370
rect 10290 4340 10440 4370
rect 10470 4340 10620 4370
rect 10650 4340 10800 4370
rect 10830 4340 10980 4370
rect 11010 4340 11160 4370
rect 11190 4340 11340 4370
rect 11370 4340 11520 4370
rect 11550 4340 11700 4370
rect 11730 4340 11880 4370
rect 11910 4340 12060 4370
rect 12090 4340 12240 4370
rect 12270 4340 12420 4370
rect 12450 4340 12600 4370
rect 12630 4340 12780 4370
rect 12810 4340 12960 4370
rect 12990 4340 13140 4370
rect 13170 4340 13320 4370
rect 13350 4340 13500 4370
rect 13530 4340 13680 4370
rect 13710 4340 13860 4370
rect 13890 4340 14040 4370
rect 14070 4340 14220 4370
rect 14250 4340 14400 4370
rect 14430 4340 14580 4370
rect 14610 4340 14760 4370
rect 14790 4340 14940 4370
rect 14970 4340 15120 4370
rect 15150 4340 15300 4370
rect 15330 4340 15480 4370
rect 15510 4340 15660 4370
rect 15690 4340 15840 4370
rect 15870 4340 16020 4370
rect 16050 4340 16200 4370
rect 16230 4340 16380 4370
rect 16410 4340 16560 4370
rect 16590 4340 16740 4370
rect 16770 4340 16920 4370
rect 16950 4340 17100 4370
rect 17130 4340 17280 4370
rect 17310 4340 17460 4370
rect 17490 4340 17640 4370
rect 17670 4340 17820 4370
rect 17850 4340 18000 4370
rect 18030 4340 18180 4370
rect 18210 4340 18360 4370
rect 18390 4340 18540 4370
rect 18570 4340 18720 4370
rect 18750 4340 18900 4370
rect 18930 4340 19080 4370
rect 19110 4340 19260 4370
rect 19290 4340 19440 4370
rect 19470 4340 19620 4370
rect 19650 4340 19800 4370
rect 19830 4340 19980 4370
rect 20010 4340 20700 4370
rect 20730 4340 20740 4370
rect 9175 4335 20740 4340
rect 9040 3450 20870 3455
rect 9040 3420 9045 3450
rect 9075 3420 9180 3450
rect 9210 3420 9900 3450
rect 9930 3420 10080 3450
rect 10110 3420 10260 3450
rect 10290 3420 10440 3450
rect 10470 3420 10620 3450
rect 10650 3420 10800 3450
rect 10830 3420 10980 3450
rect 11010 3420 11160 3450
rect 11190 3420 11340 3450
rect 11370 3420 11520 3450
rect 11550 3420 11700 3450
rect 11730 3420 11880 3450
rect 11910 3420 12060 3450
rect 12090 3420 12240 3450
rect 12270 3420 12420 3450
rect 12450 3420 12600 3450
rect 12630 3420 12780 3450
rect 12810 3420 12960 3450
rect 12990 3420 13140 3450
rect 13170 3420 13320 3450
rect 13350 3420 13500 3450
rect 13530 3420 13680 3450
rect 13710 3420 13860 3450
rect 13890 3420 14040 3450
rect 14070 3420 14220 3450
rect 14250 3420 14400 3450
rect 14430 3420 14580 3450
rect 14610 3420 14760 3450
rect 14790 3420 14940 3450
rect 14970 3420 15120 3450
rect 15150 3420 15300 3450
rect 15330 3420 15480 3450
rect 15510 3420 15660 3450
rect 15690 3420 15840 3450
rect 15870 3420 16020 3450
rect 16050 3420 16200 3450
rect 16230 3420 16380 3450
rect 16410 3420 16560 3450
rect 16590 3420 16740 3450
rect 16770 3420 16920 3450
rect 16950 3420 17100 3450
rect 17130 3420 17280 3450
rect 17310 3420 17460 3450
rect 17490 3420 17640 3450
rect 17670 3420 17820 3450
rect 17850 3420 18000 3450
rect 18030 3420 18180 3450
rect 18210 3420 18360 3450
rect 18390 3420 18540 3450
rect 18570 3420 18720 3450
rect 18750 3420 18900 3450
rect 18930 3420 19080 3450
rect 19110 3420 19260 3450
rect 19290 3420 19440 3450
rect 19470 3420 19620 3450
rect 19650 3420 19800 3450
rect 19830 3420 19980 3450
rect 20010 3420 20700 3450
rect 20730 3420 20835 3450
rect 20865 3420 20870 3450
rect 9040 3415 20870 3420
<< labels >>
rlabel locali 9185 3815 9185 3815 1 xn
rlabel locali 9185 3935 9185 3935 1 xp
rlabel locali 9185 4095 9185 4095 1 n3
rlabel locali 9185 3775 9185 3775 1 p3
rlabel locali 9185 3895 9185 3895 1 out
port 8 n
rlabel locali 9185 3735 9185 3735 1 n2
port 5 n
rlabel locali 9185 3695 9185 3695 1 n1
port 6 n
rlabel locali 9185 4015 9185 4015 1 p1
port 3 n
rlabel locali 9185 3975 9185 3975 1 p2
port 4 n
rlabel locali 9185 3855 9185 3855 1 in
port 7 n
rlabel metal2 9180 4355 9180 4355 1 VDDA
port 1 n
rlabel metal2 9180 3435 9180 3435 1 VSSA
port 2 n
<< end >>
