magic
tech sky130A
timestamp 1624035941
<< nwell >>
rect 9085 4105 20785 4385
<< mvnmos >>
rect 9195 3475 9245 3575
rect 9285 3475 9335 3575
rect 9375 3475 9425 3575
rect 9465 3475 9515 3575
rect 9555 3475 9605 3575
rect 9645 3475 9695 3575
rect 9735 3475 9785 3575
rect 9825 3475 9875 3575
rect 9915 3475 9965 3575
rect 10005 3475 10055 3575
rect 10095 3475 10145 3575
rect 10185 3475 10235 3575
rect 10275 3475 10325 3575
rect 10365 3475 10415 3575
rect 10455 3475 10505 3575
rect 10545 3475 10595 3575
rect 10635 3475 10685 3575
rect 10725 3475 10775 3575
rect 10815 3475 10865 3575
rect 10905 3475 10955 3575
rect 10995 3475 11045 3575
rect 11085 3475 11135 3575
rect 11175 3475 11225 3575
rect 11265 3475 11315 3575
rect 11355 3475 11405 3575
rect 11445 3475 11495 3575
rect 11535 3475 11585 3575
rect 11625 3475 11675 3575
rect 11715 3475 11765 3575
rect 11805 3475 11855 3575
rect 11895 3475 11945 3575
rect 11985 3475 12035 3575
rect 12075 3475 12125 3575
rect 12165 3475 12215 3575
rect 12255 3475 12305 3575
rect 12345 3475 12395 3575
rect 12435 3475 12485 3575
rect 12525 3475 12575 3575
rect 12615 3475 12665 3575
rect 12705 3475 12755 3575
rect 12795 3475 12845 3575
rect 12885 3475 12935 3575
rect 12975 3475 13025 3575
rect 13065 3475 13115 3575
rect 13155 3475 13205 3575
rect 13245 3475 13295 3575
rect 13335 3475 13385 3575
rect 13425 3475 13475 3575
rect 13515 3475 13565 3575
rect 13605 3475 13655 3575
rect 13695 3475 13745 3575
rect 13785 3475 13835 3575
rect 13875 3475 13925 3575
rect 13965 3475 14015 3575
rect 14055 3475 14105 3575
rect 14145 3475 14195 3575
rect 14235 3475 14285 3575
rect 14325 3475 14375 3575
rect 14415 3475 14465 3575
rect 14505 3475 14555 3575
rect 14595 3475 14645 3575
rect 14685 3475 14735 3575
rect 14775 3475 14825 3575
rect 14865 3475 14915 3575
rect 14955 3475 15005 3575
rect 15045 3475 15095 3575
rect 15135 3475 15185 3575
rect 15225 3475 15275 3575
rect 15315 3475 15365 3575
rect 15405 3475 15455 3575
rect 15495 3475 15545 3575
rect 15585 3475 15635 3575
rect 15675 3475 15725 3575
rect 15765 3475 15815 3575
rect 15855 3475 15905 3575
rect 15945 3475 15995 3575
rect 16035 3475 16085 3575
rect 16125 3475 16175 3575
rect 16215 3475 16265 3575
rect 16305 3475 16355 3575
rect 16395 3475 16445 3575
rect 16485 3475 16535 3575
rect 16575 3475 16625 3575
rect 16665 3475 16715 3575
rect 16755 3475 16805 3575
rect 16845 3475 16895 3575
rect 16935 3475 16985 3575
rect 17025 3475 17075 3575
rect 17115 3475 17165 3575
rect 17205 3475 17255 3575
rect 17295 3475 17345 3575
rect 17385 3475 17435 3575
rect 17475 3475 17525 3575
rect 17565 3475 17615 3575
rect 17655 3475 17705 3575
rect 17745 3475 17795 3575
rect 17835 3475 17885 3575
rect 17925 3475 17975 3575
rect 18015 3475 18065 3575
rect 18105 3475 18155 3575
rect 18195 3475 18245 3575
rect 18285 3475 18335 3575
rect 18375 3475 18425 3575
rect 18465 3475 18515 3575
rect 18555 3475 18605 3575
rect 18645 3475 18695 3575
rect 18735 3475 18785 3575
rect 18825 3475 18875 3575
rect 18915 3475 18965 3575
rect 19005 3475 19055 3575
rect 19095 3475 19145 3575
rect 19185 3475 19235 3575
rect 19275 3475 19325 3575
rect 19365 3475 19415 3575
rect 19455 3475 19505 3575
rect 19545 3475 19595 3575
rect 19635 3475 19685 3575
rect 19725 3475 19775 3575
rect 19815 3475 19865 3575
rect 19905 3475 19955 3575
rect 19995 3475 20045 3575
rect 20085 3475 20135 3575
rect 20175 3475 20225 3575
rect 20265 3475 20315 3575
rect 20355 3475 20405 3575
rect 20445 3475 20495 3575
rect 20535 3475 20585 3575
rect 20625 3475 20675 3575
<< mvpmos >>
rect 9195 4215 9245 4315
rect 9285 4215 9335 4315
rect 9375 4215 9425 4315
rect 9465 4215 9515 4315
rect 9555 4215 9605 4315
rect 9645 4215 9695 4315
rect 9735 4215 9785 4315
rect 9825 4215 9875 4315
rect 9915 4215 9965 4315
rect 10005 4215 10055 4315
rect 10095 4215 10145 4315
rect 10185 4215 10235 4315
rect 10275 4215 10325 4315
rect 10365 4215 10415 4315
rect 10455 4215 10505 4315
rect 10545 4215 10595 4315
rect 10635 4215 10685 4315
rect 10725 4215 10775 4315
rect 10815 4215 10865 4315
rect 10905 4215 10955 4315
rect 10995 4215 11045 4315
rect 11085 4215 11135 4315
rect 11175 4215 11225 4315
rect 11265 4215 11315 4315
rect 11355 4215 11405 4315
rect 11445 4215 11495 4315
rect 11535 4215 11585 4315
rect 11625 4215 11675 4315
rect 11715 4215 11765 4315
rect 11805 4215 11855 4315
rect 11895 4215 11945 4315
rect 11985 4215 12035 4315
rect 12075 4215 12125 4315
rect 12165 4215 12215 4315
rect 12255 4215 12305 4315
rect 12345 4215 12395 4315
rect 12435 4215 12485 4315
rect 12525 4215 12575 4315
rect 12615 4215 12665 4315
rect 12705 4215 12755 4315
rect 12795 4215 12845 4315
rect 12885 4215 12935 4315
rect 12975 4215 13025 4315
rect 13065 4215 13115 4315
rect 13155 4215 13205 4315
rect 13245 4215 13295 4315
rect 13335 4215 13385 4315
rect 13425 4215 13475 4315
rect 13515 4215 13565 4315
rect 13605 4215 13655 4315
rect 13695 4215 13745 4315
rect 13785 4215 13835 4315
rect 13875 4215 13925 4315
rect 13965 4215 14015 4315
rect 14055 4215 14105 4315
rect 14145 4215 14195 4315
rect 14235 4215 14285 4315
rect 14325 4215 14375 4315
rect 14415 4215 14465 4315
rect 14505 4215 14555 4315
rect 14595 4215 14645 4315
rect 14685 4215 14735 4315
rect 14775 4215 14825 4315
rect 14865 4215 14915 4315
rect 14955 4215 15005 4315
rect 15045 4215 15095 4315
rect 15135 4215 15185 4315
rect 15225 4215 15275 4315
rect 15315 4215 15365 4315
rect 15405 4215 15455 4315
rect 15495 4215 15545 4315
rect 15585 4215 15635 4315
rect 15675 4215 15725 4315
rect 15765 4215 15815 4315
rect 15855 4215 15905 4315
rect 15945 4215 15995 4315
rect 16035 4215 16085 4315
rect 16125 4215 16175 4315
rect 16215 4215 16265 4315
rect 16305 4215 16355 4315
rect 16395 4215 16445 4315
rect 16485 4215 16535 4315
rect 16575 4215 16625 4315
rect 16665 4215 16715 4315
rect 16755 4215 16805 4315
rect 16845 4215 16895 4315
rect 16935 4215 16985 4315
rect 17025 4215 17075 4315
rect 17115 4215 17165 4315
rect 17205 4215 17255 4315
rect 17295 4215 17345 4315
rect 17385 4215 17435 4315
rect 17475 4215 17525 4315
rect 17565 4215 17615 4315
rect 17655 4215 17705 4315
rect 17745 4215 17795 4315
rect 17835 4215 17885 4315
rect 17925 4215 17975 4315
rect 18015 4215 18065 4315
rect 18105 4215 18155 4315
rect 18195 4215 18245 4315
rect 18285 4215 18335 4315
rect 18375 4215 18425 4315
rect 18465 4215 18515 4315
rect 18555 4215 18605 4315
rect 18645 4215 18695 4315
rect 18735 4215 18785 4315
rect 18825 4215 18875 4315
rect 18915 4215 18965 4315
rect 19005 4215 19055 4315
rect 19095 4215 19145 4315
rect 19185 4215 19235 4315
rect 19275 4215 19325 4315
rect 19365 4215 19415 4315
rect 19455 4215 19505 4315
rect 19545 4215 19595 4315
rect 19635 4215 19685 4315
rect 19725 4215 19775 4315
rect 19815 4215 19865 4315
rect 19905 4215 19955 4315
rect 19995 4215 20045 4315
rect 20085 4215 20135 4315
rect 20175 4215 20225 4315
rect 20265 4215 20315 4315
rect 20355 4215 20405 4315
rect 20445 4215 20495 4315
rect 20535 4215 20585 4315
rect 20625 4215 20675 4315
<< mvndiff >>
rect 9155 3565 9195 3575
rect 9155 3485 9165 3565
rect 9185 3485 9195 3565
rect 9155 3475 9195 3485
rect 9245 3565 9285 3575
rect 9245 3485 9255 3565
rect 9275 3485 9285 3565
rect 9245 3475 9285 3485
rect 9335 3565 9375 3575
rect 9335 3485 9345 3565
rect 9365 3485 9375 3565
rect 9335 3475 9375 3485
rect 9425 3565 9465 3575
rect 9425 3485 9435 3565
rect 9455 3485 9465 3565
rect 9425 3475 9465 3485
rect 9515 3565 9555 3575
rect 9515 3485 9525 3565
rect 9545 3485 9555 3565
rect 9515 3475 9555 3485
rect 9605 3565 9645 3575
rect 9605 3485 9615 3565
rect 9635 3485 9645 3565
rect 9605 3475 9645 3485
rect 9695 3565 9735 3575
rect 9695 3485 9705 3565
rect 9725 3485 9735 3565
rect 9695 3475 9735 3485
rect 9785 3565 9825 3575
rect 9785 3485 9795 3565
rect 9815 3485 9825 3565
rect 9785 3475 9825 3485
rect 9875 3565 9915 3575
rect 9875 3485 9885 3565
rect 9905 3485 9915 3565
rect 9875 3475 9915 3485
rect 9965 3565 10005 3575
rect 9965 3485 9975 3565
rect 9995 3485 10005 3565
rect 9965 3475 10005 3485
rect 10055 3565 10095 3575
rect 10055 3485 10065 3565
rect 10085 3485 10095 3565
rect 10055 3475 10095 3485
rect 10145 3565 10185 3575
rect 10145 3485 10155 3565
rect 10175 3485 10185 3565
rect 10145 3475 10185 3485
rect 10235 3565 10275 3575
rect 10235 3485 10245 3565
rect 10265 3485 10275 3565
rect 10235 3475 10275 3485
rect 10325 3565 10365 3575
rect 10325 3485 10335 3565
rect 10355 3485 10365 3565
rect 10325 3475 10365 3485
rect 10415 3565 10455 3575
rect 10415 3485 10425 3565
rect 10445 3485 10455 3565
rect 10415 3475 10455 3485
rect 10505 3565 10545 3575
rect 10505 3485 10515 3565
rect 10535 3485 10545 3565
rect 10505 3475 10545 3485
rect 10595 3565 10635 3575
rect 10595 3485 10605 3565
rect 10625 3485 10635 3565
rect 10595 3475 10635 3485
rect 10685 3565 10725 3575
rect 10685 3485 10695 3565
rect 10715 3485 10725 3565
rect 10685 3475 10725 3485
rect 10775 3565 10815 3575
rect 10775 3485 10785 3565
rect 10805 3485 10815 3565
rect 10775 3475 10815 3485
rect 10865 3565 10905 3575
rect 10865 3485 10875 3565
rect 10895 3485 10905 3565
rect 10865 3475 10905 3485
rect 10955 3565 10995 3575
rect 10955 3485 10965 3565
rect 10985 3485 10995 3565
rect 10955 3475 10995 3485
rect 11045 3565 11085 3575
rect 11045 3485 11055 3565
rect 11075 3485 11085 3565
rect 11045 3475 11085 3485
rect 11135 3565 11175 3575
rect 11135 3485 11145 3565
rect 11165 3485 11175 3565
rect 11135 3475 11175 3485
rect 11225 3565 11265 3575
rect 11225 3485 11235 3565
rect 11255 3485 11265 3565
rect 11225 3475 11265 3485
rect 11315 3565 11355 3575
rect 11315 3485 11325 3565
rect 11345 3485 11355 3565
rect 11315 3475 11355 3485
rect 11405 3565 11445 3575
rect 11405 3485 11415 3565
rect 11435 3485 11445 3565
rect 11405 3475 11445 3485
rect 11495 3565 11535 3575
rect 11495 3485 11505 3565
rect 11525 3485 11535 3565
rect 11495 3475 11535 3485
rect 11585 3565 11625 3575
rect 11585 3485 11595 3565
rect 11615 3485 11625 3565
rect 11585 3475 11625 3485
rect 11675 3565 11715 3575
rect 11675 3485 11685 3565
rect 11705 3485 11715 3565
rect 11675 3475 11715 3485
rect 11765 3565 11805 3575
rect 11765 3485 11775 3565
rect 11795 3485 11805 3565
rect 11765 3475 11805 3485
rect 11855 3565 11895 3575
rect 11855 3485 11865 3565
rect 11885 3485 11895 3565
rect 11855 3475 11895 3485
rect 11945 3565 11985 3575
rect 11945 3485 11955 3565
rect 11975 3485 11985 3565
rect 11945 3475 11985 3485
rect 12035 3565 12075 3575
rect 12035 3485 12045 3565
rect 12065 3485 12075 3565
rect 12035 3475 12075 3485
rect 12125 3565 12165 3575
rect 12125 3485 12135 3565
rect 12155 3485 12165 3565
rect 12125 3475 12165 3485
rect 12215 3565 12255 3575
rect 12215 3485 12225 3565
rect 12245 3485 12255 3565
rect 12215 3475 12255 3485
rect 12305 3565 12345 3575
rect 12305 3485 12315 3565
rect 12335 3485 12345 3565
rect 12305 3475 12345 3485
rect 12395 3565 12435 3575
rect 12395 3485 12405 3565
rect 12425 3485 12435 3565
rect 12395 3475 12435 3485
rect 12485 3565 12525 3575
rect 12485 3485 12495 3565
rect 12515 3485 12525 3565
rect 12485 3475 12525 3485
rect 12575 3565 12615 3575
rect 12575 3485 12585 3565
rect 12605 3485 12615 3565
rect 12575 3475 12615 3485
rect 12665 3565 12705 3575
rect 12665 3485 12675 3565
rect 12695 3485 12705 3565
rect 12665 3475 12705 3485
rect 12755 3565 12795 3575
rect 12755 3485 12765 3565
rect 12785 3485 12795 3565
rect 12755 3475 12795 3485
rect 12845 3565 12885 3575
rect 12845 3485 12855 3565
rect 12875 3485 12885 3565
rect 12845 3475 12885 3485
rect 12935 3565 12975 3575
rect 12935 3485 12945 3565
rect 12965 3485 12975 3565
rect 12935 3475 12975 3485
rect 13025 3565 13065 3575
rect 13025 3485 13035 3565
rect 13055 3485 13065 3565
rect 13025 3475 13065 3485
rect 13115 3565 13155 3575
rect 13115 3485 13125 3565
rect 13145 3485 13155 3565
rect 13115 3475 13155 3485
rect 13205 3565 13245 3575
rect 13205 3485 13215 3565
rect 13235 3485 13245 3565
rect 13205 3475 13245 3485
rect 13295 3565 13335 3575
rect 13295 3485 13305 3565
rect 13325 3485 13335 3565
rect 13295 3475 13335 3485
rect 13385 3565 13425 3575
rect 13385 3485 13395 3565
rect 13415 3485 13425 3565
rect 13385 3475 13425 3485
rect 13475 3565 13515 3575
rect 13475 3485 13485 3565
rect 13505 3485 13515 3565
rect 13475 3475 13515 3485
rect 13565 3565 13605 3575
rect 13565 3485 13575 3565
rect 13595 3485 13605 3565
rect 13565 3475 13605 3485
rect 13655 3565 13695 3575
rect 13655 3485 13665 3565
rect 13685 3485 13695 3565
rect 13655 3475 13695 3485
rect 13745 3565 13785 3575
rect 13745 3485 13755 3565
rect 13775 3485 13785 3565
rect 13745 3475 13785 3485
rect 13835 3565 13875 3575
rect 13835 3485 13845 3565
rect 13865 3485 13875 3565
rect 13835 3475 13875 3485
rect 13925 3565 13965 3575
rect 13925 3485 13935 3565
rect 13955 3485 13965 3565
rect 13925 3475 13965 3485
rect 14015 3565 14055 3575
rect 14015 3485 14025 3565
rect 14045 3485 14055 3565
rect 14015 3475 14055 3485
rect 14105 3565 14145 3575
rect 14105 3485 14115 3565
rect 14135 3485 14145 3565
rect 14105 3475 14145 3485
rect 14195 3565 14235 3575
rect 14195 3485 14205 3565
rect 14225 3485 14235 3565
rect 14195 3475 14235 3485
rect 14285 3565 14325 3575
rect 14285 3485 14295 3565
rect 14315 3485 14325 3565
rect 14285 3475 14325 3485
rect 14375 3565 14415 3575
rect 14375 3485 14385 3565
rect 14405 3485 14415 3565
rect 14375 3475 14415 3485
rect 14465 3565 14505 3575
rect 14465 3485 14475 3565
rect 14495 3485 14505 3565
rect 14465 3475 14505 3485
rect 14555 3565 14595 3575
rect 14555 3485 14565 3565
rect 14585 3485 14595 3565
rect 14555 3475 14595 3485
rect 14645 3565 14685 3575
rect 14645 3485 14655 3565
rect 14675 3485 14685 3565
rect 14645 3475 14685 3485
rect 14735 3565 14775 3575
rect 14735 3485 14745 3565
rect 14765 3485 14775 3565
rect 14735 3475 14775 3485
rect 14825 3565 14865 3575
rect 14825 3485 14835 3565
rect 14855 3485 14865 3565
rect 14825 3475 14865 3485
rect 14915 3565 14955 3575
rect 14915 3485 14925 3565
rect 14945 3485 14955 3565
rect 14915 3475 14955 3485
rect 15005 3565 15045 3575
rect 15005 3485 15015 3565
rect 15035 3485 15045 3565
rect 15005 3475 15045 3485
rect 15095 3565 15135 3575
rect 15095 3485 15105 3565
rect 15125 3485 15135 3565
rect 15095 3475 15135 3485
rect 15185 3565 15225 3575
rect 15185 3485 15195 3565
rect 15215 3485 15225 3565
rect 15185 3475 15225 3485
rect 15275 3565 15315 3575
rect 15275 3485 15285 3565
rect 15305 3485 15315 3565
rect 15275 3475 15315 3485
rect 15365 3565 15405 3575
rect 15365 3485 15375 3565
rect 15395 3485 15405 3565
rect 15365 3475 15405 3485
rect 15455 3565 15495 3575
rect 15455 3485 15465 3565
rect 15485 3485 15495 3565
rect 15455 3475 15495 3485
rect 15545 3565 15585 3575
rect 15545 3485 15555 3565
rect 15575 3485 15585 3565
rect 15545 3475 15585 3485
rect 15635 3565 15675 3575
rect 15635 3485 15645 3565
rect 15665 3485 15675 3565
rect 15635 3475 15675 3485
rect 15725 3565 15765 3575
rect 15725 3485 15735 3565
rect 15755 3485 15765 3565
rect 15725 3475 15765 3485
rect 15815 3565 15855 3575
rect 15815 3485 15825 3565
rect 15845 3485 15855 3565
rect 15815 3475 15855 3485
rect 15905 3565 15945 3575
rect 15905 3485 15915 3565
rect 15935 3485 15945 3565
rect 15905 3475 15945 3485
rect 15995 3565 16035 3575
rect 15995 3485 16005 3565
rect 16025 3485 16035 3565
rect 15995 3475 16035 3485
rect 16085 3565 16125 3575
rect 16085 3485 16095 3565
rect 16115 3485 16125 3565
rect 16085 3475 16125 3485
rect 16175 3565 16215 3575
rect 16175 3485 16185 3565
rect 16205 3485 16215 3565
rect 16175 3475 16215 3485
rect 16265 3565 16305 3575
rect 16265 3485 16275 3565
rect 16295 3485 16305 3565
rect 16265 3475 16305 3485
rect 16355 3565 16395 3575
rect 16355 3485 16365 3565
rect 16385 3485 16395 3565
rect 16355 3475 16395 3485
rect 16445 3565 16485 3575
rect 16445 3485 16455 3565
rect 16475 3485 16485 3565
rect 16445 3475 16485 3485
rect 16535 3565 16575 3575
rect 16535 3485 16545 3565
rect 16565 3485 16575 3565
rect 16535 3475 16575 3485
rect 16625 3565 16665 3575
rect 16625 3485 16635 3565
rect 16655 3485 16665 3565
rect 16625 3475 16665 3485
rect 16715 3565 16755 3575
rect 16715 3485 16725 3565
rect 16745 3485 16755 3565
rect 16715 3475 16755 3485
rect 16805 3565 16845 3575
rect 16805 3485 16815 3565
rect 16835 3485 16845 3565
rect 16805 3475 16845 3485
rect 16895 3565 16935 3575
rect 16895 3485 16905 3565
rect 16925 3485 16935 3565
rect 16895 3475 16935 3485
rect 16985 3565 17025 3575
rect 16985 3485 16995 3565
rect 17015 3485 17025 3565
rect 16985 3475 17025 3485
rect 17075 3565 17115 3575
rect 17075 3485 17085 3565
rect 17105 3485 17115 3565
rect 17075 3475 17115 3485
rect 17165 3565 17205 3575
rect 17165 3485 17175 3565
rect 17195 3485 17205 3565
rect 17165 3475 17205 3485
rect 17255 3565 17295 3575
rect 17255 3485 17265 3565
rect 17285 3485 17295 3565
rect 17255 3475 17295 3485
rect 17345 3565 17385 3575
rect 17345 3485 17355 3565
rect 17375 3485 17385 3565
rect 17345 3475 17385 3485
rect 17435 3565 17475 3575
rect 17435 3485 17445 3565
rect 17465 3485 17475 3565
rect 17435 3475 17475 3485
rect 17525 3565 17565 3575
rect 17525 3485 17535 3565
rect 17555 3485 17565 3565
rect 17525 3475 17565 3485
rect 17615 3565 17655 3575
rect 17615 3485 17625 3565
rect 17645 3485 17655 3565
rect 17615 3475 17655 3485
rect 17705 3565 17745 3575
rect 17705 3485 17715 3565
rect 17735 3485 17745 3565
rect 17705 3475 17745 3485
rect 17795 3565 17835 3575
rect 17795 3485 17805 3565
rect 17825 3485 17835 3565
rect 17795 3475 17835 3485
rect 17885 3565 17925 3575
rect 17885 3485 17895 3565
rect 17915 3485 17925 3565
rect 17885 3475 17925 3485
rect 17975 3565 18015 3575
rect 17975 3485 17985 3565
rect 18005 3485 18015 3565
rect 17975 3475 18015 3485
rect 18065 3565 18105 3575
rect 18065 3485 18075 3565
rect 18095 3485 18105 3565
rect 18065 3475 18105 3485
rect 18155 3565 18195 3575
rect 18155 3485 18165 3565
rect 18185 3485 18195 3565
rect 18155 3475 18195 3485
rect 18245 3565 18285 3575
rect 18245 3485 18255 3565
rect 18275 3485 18285 3565
rect 18245 3475 18285 3485
rect 18335 3565 18375 3575
rect 18335 3485 18345 3565
rect 18365 3485 18375 3565
rect 18335 3475 18375 3485
rect 18425 3565 18465 3575
rect 18425 3485 18435 3565
rect 18455 3485 18465 3565
rect 18425 3475 18465 3485
rect 18515 3565 18555 3575
rect 18515 3485 18525 3565
rect 18545 3485 18555 3565
rect 18515 3475 18555 3485
rect 18605 3565 18645 3575
rect 18605 3485 18615 3565
rect 18635 3485 18645 3565
rect 18605 3475 18645 3485
rect 18695 3565 18735 3575
rect 18695 3485 18705 3565
rect 18725 3485 18735 3565
rect 18695 3475 18735 3485
rect 18785 3565 18825 3575
rect 18785 3485 18795 3565
rect 18815 3485 18825 3565
rect 18785 3475 18825 3485
rect 18875 3565 18915 3575
rect 18875 3485 18885 3565
rect 18905 3485 18915 3565
rect 18875 3475 18915 3485
rect 18965 3565 19005 3575
rect 18965 3485 18975 3565
rect 18995 3485 19005 3565
rect 18965 3475 19005 3485
rect 19055 3565 19095 3575
rect 19055 3485 19065 3565
rect 19085 3485 19095 3565
rect 19055 3475 19095 3485
rect 19145 3565 19185 3575
rect 19145 3485 19155 3565
rect 19175 3485 19185 3565
rect 19145 3475 19185 3485
rect 19235 3565 19275 3575
rect 19235 3485 19245 3565
rect 19265 3485 19275 3565
rect 19235 3475 19275 3485
rect 19325 3565 19365 3575
rect 19325 3485 19335 3565
rect 19355 3485 19365 3565
rect 19325 3475 19365 3485
rect 19415 3565 19455 3575
rect 19415 3485 19425 3565
rect 19445 3485 19455 3565
rect 19415 3475 19455 3485
rect 19505 3565 19545 3575
rect 19505 3485 19515 3565
rect 19535 3485 19545 3565
rect 19505 3475 19545 3485
rect 19595 3565 19635 3575
rect 19595 3485 19605 3565
rect 19625 3485 19635 3565
rect 19595 3475 19635 3485
rect 19685 3565 19725 3575
rect 19685 3485 19695 3565
rect 19715 3485 19725 3565
rect 19685 3475 19725 3485
rect 19775 3565 19815 3575
rect 19775 3485 19785 3565
rect 19805 3485 19815 3565
rect 19775 3475 19815 3485
rect 19865 3565 19905 3575
rect 19865 3485 19875 3565
rect 19895 3485 19905 3565
rect 19865 3475 19905 3485
rect 19955 3565 19995 3575
rect 19955 3485 19965 3565
rect 19985 3485 19995 3565
rect 19955 3475 19995 3485
rect 20045 3565 20085 3575
rect 20045 3485 20055 3565
rect 20075 3485 20085 3565
rect 20045 3475 20085 3485
rect 20135 3565 20175 3575
rect 20135 3485 20145 3565
rect 20165 3485 20175 3565
rect 20135 3475 20175 3485
rect 20225 3565 20265 3575
rect 20225 3485 20235 3565
rect 20255 3485 20265 3565
rect 20225 3475 20265 3485
rect 20315 3565 20355 3575
rect 20315 3485 20325 3565
rect 20345 3485 20355 3565
rect 20315 3475 20355 3485
rect 20405 3565 20445 3575
rect 20405 3485 20415 3565
rect 20435 3485 20445 3565
rect 20405 3475 20445 3485
rect 20495 3565 20535 3575
rect 20495 3485 20505 3565
rect 20525 3485 20535 3565
rect 20495 3475 20535 3485
rect 20585 3565 20625 3575
rect 20585 3485 20595 3565
rect 20615 3485 20625 3565
rect 20585 3475 20625 3485
rect 20675 3565 20715 3575
rect 20675 3485 20685 3565
rect 20705 3485 20715 3565
rect 20675 3475 20715 3485
<< mvpdiff >>
rect 9155 4305 9195 4315
rect 9155 4225 9165 4305
rect 9185 4225 9195 4305
rect 9155 4215 9195 4225
rect 9245 4305 9285 4315
rect 9245 4225 9255 4305
rect 9275 4225 9285 4305
rect 9245 4215 9285 4225
rect 9335 4305 9375 4315
rect 9335 4225 9345 4305
rect 9365 4225 9375 4305
rect 9335 4215 9375 4225
rect 9425 4305 9465 4315
rect 9425 4225 9435 4305
rect 9455 4225 9465 4305
rect 9425 4215 9465 4225
rect 9515 4305 9555 4315
rect 9515 4225 9525 4305
rect 9545 4225 9555 4305
rect 9515 4215 9555 4225
rect 9605 4305 9645 4315
rect 9605 4225 9615 4305
rect 9635 4225 9645 4305
rect 9605 4215 9645 4225
rect 9695 4305 9735 4315
rect 9695 4225 9705 4305
rect 9725 4225 9735 4305
rect 9695 4215 9735 4225
rect 9785 4305 9825 4315
rect 9785 4225 9795 4305
rect 9815 4225 9825 4305
rect 9785 4215 9825 4225
rect 9875 4305 9915 4315
rect 9875 4225 9885 4305
rect 9905 4225 9915 4305
rect 9875 4215 9915 4225
rect 9965 4305 10005 4315
rect 9965 4225 9975 4305
rect 9995 4225 10005 4305
rect 9965 4215 10005 4225
rect 10055 4305 10095 4315
rect 10055 4225 10065 4305
rect 10085 4225 10095 4305
rect 10055 4215 10095 4225
rect 10145 4305 10185 4315
rect 10145 4225 10155 4305
rect 10175 4225 10185 4305
rect 10145 4215 10185 4225
rect 10235 4305 10275 4315
rect 10235 4225 10245 4305
rect 10265 4225 10275 4305
rect 10235 4215 10275 4225
rect 10325 4305 10365 4315
rect 10325 4225 10335 4305
rect 10355 4225 10365 4305
rect 10325 4215 10365 4225
rect 10415 4305 10455 4315
rect 10415 4225 10425 4305
rect 10445 4225 10455 4305
rect 10415 4215 10455 4225
rect 10505 4305 10545 4315
rect 10505 4225 10515 4305
rect 10535 4225 10545 4305
rect 10505 4215 10545 4225
rect 10595 4305 10635 4315
rect 10595 4225 10605 4305
rect 10625 4225 10635 4305
rect 10595 4215 10635 4225
rect 10685 4305 10725 4315
rect 10685 4225 10695 4305
rect 10715 4225 10725 4305
rect 10685 4215 10725 4225
rect 10775 4305 10815 4315
rect 10775 4225 10785 4305
rect 10805 4225 10815 4305
rect 10775 4215 10815 4225
rect 10865 4305 10905 4315
rect 10865 4225 10875 4305
rect 10895 4225 10905 4305
rect 10865 4215 10905 4225
rect 10955 4305 10995 4315
rect 10955 4225 10965 4305
rect 10985 4225 10995 4305
rect 10955 4215 10995 4225
rect 11045 4305 11085 4315
rect 11045 4225 11055 4305
rect 11075 4225 11085 4305
rect 11045 4215 11085 4225
rect 11135 4305 11175 4315
rect 11135 4225 11145 4305
rect 11165 4225 11175 4305
rect 11135 4215 11175 4225
rect 11225 4305 11265 4315
rect 11225 4225 11235 4305
rect 11255 4225 11265 4305
rect 11225 4215 11265 4225
rect 11315 4305 11355 4315
rect 11315 4225 11325 4305
rect 11345 4225 11355 4305
rect 11315 4215 11355 4225
rect 11405 4305 11445 4315
rect 11405 4225 11415 4305
rect 11435 4225 11445 4305
rect 11405 4215 11445 4225
rect 11495 4305 11535 4315
rect 11495 4225 11505 4305
rect 11525 4225 11535 4305
rect 11495 4215 11535 4225
rect 11585 4305 11625 4315
rect 11585 4225 11595 4305
rect 11615 4225 11625 4305
rect 11585 4215 11625 4225
rect 11675 4305 11715 4315
rect 11675 4225 11685 4305
rect 11705 4225 11715 4305
rect 11675 4215 11715 4225
rect 11765 4305 11805 4315
rect 11765 4225 11775 4305
rect 11795 4225 11805 4305
rect 11765 4215 11805 4225
rect 11855 4305 11895 4315
rect 11855 4225 11865 4305
rect 11885 4225 11895 4305
rect 11855 4215 11895 4225
rect 11945 4305 11985 4315
rect 11945 4225 11955 4305
rect 11975 4225 11985 4305
rect 11945 4215 11985 4225
rect 12035 4305 12075 4315
rect 12035 4225 12045 4305
rect 12065 4225 12075 4305
rect 12035 4215 12075 4225
rect 12125 4305 12165 4315
rect 12125 4225 12135 4305
rect 12155 4225 12165 4305
rect 12125 4215 12165 4225
rect 12215 4305 12255 4315
rect 12215 4225 12225 4305
rect 12245 4225 12255 4305
rect 12215 4215 12255 4225
rect 12305 4305 12345 4315
rect 12305 4225 12315 4305
rect 12335 4225 12345 4305
rect 12305 4215 12345 4225
rect 12395 4305 12435 4315
rect 12395 4225 12405 4305
rect 12425 4225 12435 4305
rect 12395 4215 12435 4225
rect 12485 4305 12525 4315
rect 12485 4225 12495 4305
rect 12515 4225 12525 4305
rect 12485 4215 12525 4225
rect 12575 4305 12615 4315
rect 12575 4225 12585 4305
rect 12605 4225 12615 4305
rect 12575 4215 12615 4225
rect 12665 4305 12705 4315
rect 12665 4225 12675 4305
rect 12695 4225 12705 4305
rect 12665 4215 12705 4225
rect 12755 4305 12795 4315
rect 12755 4225 12765 4305
rect 12785 4225 12795 4305
rect 12755 4215 12795 4225
rect 12845 4305 12885 4315
rect 12845 4225 12855 4305
rect 12875 4225 12885 4305
rect 12845 4215 12885 4225
rect 12935 4305 12975 4315
rect 12935 4225 12945 4305
rect 12965 4225 12975 4305
rect 12935 4215 12975 4225
rect 13025 4305 13065 4315
rect 13025 4225 13035 4305
rect 13055 4225 13065 4305
rect 13025 4215 13065 4225
rect 13115 4305 13155 4315
rect 13115 4225 13125 4305
rect 13145 4225 13155 4305
rect 13115 4215 13155 4225
rect 13205 4305 13245 4315
rect 13205 4225 13215 4305
rect 13235 4225 13245 4305
rect 13205 4215 13245 4225
rect 13295 4305 13335 4315
rect 13295 4225 13305 4305
rect 13325 4225 13335 4305
rect 13295 4215 13335 4225
rect 13385 4305 13425 4315
rect 13385 4225 13395 4305
rect 13415 4225 13425 4305
rect 13385 4215 13425 4225
rect 13475 4305 13515 4315
rect 13475 4225 13485 4305
rect 13505 4225 13515 4305
rect 13475 4215 13515 4225
rect 13565 4305 13605 4315
rect 13565 4225 13575 4305
rect 13595 4225 13605 4305
rect 13565 4215 13605 4225
rect 13655 4305 13695 4315
rect 13655 4225 13665 4305
rect 13685 4225 13695 4305
rect 13655 4215 13695 4225
rect 13745 4305 13785 4315
rect 13745 4225 13755 4305
rect 13775 4225 13785 4305
rect 13745 4215 13785 4225
rect 13835 4305 13875 4315
rect 13835 4225 13845 4305
rect 13865 4225 13875 4305
rect 13835 4215 13875 4225
rect 13925 4305 13965 4315
rect 13925 4225 13935 4305
rect 13955 4225 13965 4305
rect 13925 4215 13965 4225
rect 14015 4305 14055 4315
rect 14015 4225 14025 4305
rect 14045 4225 14055 4305
rect 14015 4215 14055 4225
rect 14105 4305 14145 4315
rect 14105 4225 14115 4305
rect 14135 4225 14145 4305
rect 14105 4215 14145 4225
rect 14195 4305 14235 4315
rect 14195 4225 14205 4305
rect 14225 4225 14235 4305
rect 14195 4215 14235 4225
rect 14285 4305 14325 4315
rect 14285 4225 14295 4305
rect 14315 4225 14325 4305
rect 14285 4215 14325 4225
rect 14375 4305 14415 4315
rect 14375 4225 14385 4305
rect 14405 4225 14415 4305
rect 14375 4215 14415 4225
rect 14465 4305 14505 4315
rect 14465 4225 14475 4305
rect 14495 4225 14505 4305
rect 14465 4215 14505 4225
rect 14555 4305 14595 4315
rect 14555 4225 14565 4305
rect 14585 4225 14595 4305
rect 14555 4215 14595 4225
rect 14645 4305 14685 4315
rect 14645 4225 14655 4305
rect 14675 4225 14685 4305
rect 14645 4215 14685 4225
rect 14735 4305 14775 4315
rect 14735 4225 14745 4305
rect 14765 4225 14775 4305
rect 14735 4215 14775 4225
rect 14825 4305 14865 4315
rect 14825 4225 14835 4305
rect 14855 4225 14865 4305
rect 14825 4215 14865 4225
rect 14915 4305 14955 4315
rect 14915 4225 14925 4305
rect 14945 4225 14955 4305
rect 14915 4215 14955 4225
rect 15005 4305 15045 4315
rect 15005 4225 15015 4305
rect 15035 4225 15045 4305
rect 15005 4215 15045 4225
rect 15095 4305 15135 4315
rect 15095 4225 15105 4305
rect 15125 4225 15135 4305
rect 15095 4215 15135 4225
rect 15185 4305 15225 4315
rect 15185 4225 15195 4305
rect 15215 4225 15225 4305
rect 15185 4215 15225 4225
rect 15275 4305 15315 4315
rect 15275 4225 15285 4305
rect 15305 4225 15315 4305
rect 15275 4215 15315 4225
rect 15365 4305 15405 4315
rect 15365 4225 15375 4305
rect 15395 4225 15405 4305
rect 15365 4215 15405 4225
rect 15455 4305 15495 4315
rect 15455 4225 15465 4305
rect 15485 4225 15495 4305
rect 15455 4215 15495 4225
rect 15545 4305 15585 4315
rect 15545 4225 15555 4305
rect 15575 4225 15585 4305
rect 15545 4215 15585 4225
rect 15635 4305 15675 4315
rect 15635 4225 15645 4305
rect 15665 4225 15675 4305
rect 15635 4215 15675 4225
rect 15725 4305 15765 4315
rect 15725 4225 15735 4305
rect 15755 4225 15765 4305
rect 15725 4215 15765 4225
rect 15815 4305 15855 4315
rect 15815 4225 15825 4305
rect 15845 4225 15855 4305
rect 15815 4215 15855 4225
rect 15905 4305 15945 4315
rect 15905 4225 15915 4305
rect 15935 4225 15945 4305
rect 15905 4215 15945 4225
rect 15995 4305 16035 4315
rect 15995 4225 16005 4305
rect 16025 4225 16035 4305
rect 15995 4215 16035 4225
rect 16085 4305 16125 4315
rect 16085 4225 16095 4305
rect 16115 4225 16125 4305
rect 16085 4215 16125 4225
rect 16175 4305 16215 4315
rect 16175 4225 16185 4305
rect 16205 4225 16215 4305
rect 16175 4215 16215 4225
rect 16265 4305 16305 4315
rect 16265 4225 16275 4305
rect 16295 4225 16305 4305
rect 16265 4215 16305 4225
rect 16355 4305 16395 4315
rect 16355 4225 16365 4305
rect 16385 4225 16395 4305
rect 16355 4215 16395 4225
rect 16445 4305 16485 4315
rect 16445 4225 16455 4305
rect 16475 4225 16485 4305
rect 16445 4215 16485 4225
rect 16535 4305 16575 4315
rect 16535 4225 16545 4305
rect 16565 4225 16575 4305
rect 16535 4215 16575 4225
rect 16625 4305 16665 4315
rect 16625 4225 16635 4305
rect 16655 4225 16665 4305
rect 16625 4215 16665 4225
rect 16715 4305 16755 4315
rect 16715 4225 16725 4305
rect 16745 4225 16755 4305
rect 16715 4215 16755 4225
rect 16805 4305 16845 4315
rect 16805 4225 16815 4305
rect 16835 4225 16845 4305
rect 16805 4215 16845 4225
rect 16895 4305 16935 4315
rect 16895 4225 16905 4305
rect 16925 4225 16935 4305
rect 16895 4215 16935 4225
rect 16985 4305 17025 4315
rect 16985 4225 16995 4305
rect 17015 4225 17025 4305
rect 16985 4215 17025 4225
rect 17075 4305 17115 4315
rect 17075 4225 17085 4305
rect 17105 4225 17115 4305
rect 17075 4215 17115 4225
rect 17165 4305 17205 4315
rect 17165 4225 17175 4305
rect 17195 4225 17205 4305
rect 17165 4215 17205 4225
rect 17255 4305 17295 4315
rect 17255 4225 17265 4305
rect 17285 4225 17295 4305
rect 17255 4215 17295 4225
rect 17345 4305 17385 4315
rect 17345 4225 17355 4305
rect 17375 4225 17385 4305
rect 17345 4215 17385 4225
rect 17435 4305 17475 4315
rect 17435 4225 17445 4305
rect 17465 4225 17475 4305
rect 17435 4215 17475 4225
rect 17525 4305 17565 4315
rect 17525 4225 17535 4305
rect 17555 4225 17565 4305
rect 17525 4215 17565 4225
rect 17615 4305 17655 4315
rect 17615 4225 17625 4305
rect 17645 4225 17655 4305
rect 17615 4215 17655 4225
rect 17705 4305 17745 4315
rect 17705 4225 17715 4305
rect 17735 4225 17745 4305
rect 17705 4215 17745 4225
rect 17795 4305 17835 4315
rect 17795 4225 17805 4305
rect 17825 4225 17835 4305
rect 17795 4215 17835 4225
rect 17885 4305 17925 4315
rect 17885 4225 17895 4305
rect 17915 4225 17925 4305
rect 17885 4215 17925 4225
rect 17975 4305 18015 4315
rect 17975 4225 17985 4305
rect 18005 4225 18015 4305
rect 17975 4215 18015 4225
rect 18065 4305 18105 4315
rect 18065 4225 18075 4305
rect 18095 4225 18105 4305
rect 18065 4215 18105 4225
rect 18155 4305 18195 4315
rect 18155 4225 18165 4305
rect 18185 4225 18195 4305
rect 18155 4215 18195 4225
rect 18245 4305 18285 4315
rect 18245 4225 18255 4305
rect 18275 4225 18285 4305
rect 18245 4215 18285 4225
rect 18335 4305 18375 4315
rect 18335 4225 18345 4305
rect 18365 4225 18375 4305
rect 18335 4215 18375 4225
rect 18425 4305 18465 4315
rect 18425 4225 18435 4305
rect 18455 4225 18465 4305
rect 18425 4215 18465 4225
rect 18515 4305 18555 4315
rect 18515 4225 18525 4305
rect 18545 4225 18555 4305
rect 18515 4215 18555 4225
rect 18605 4305 18645 4315
rect 18605 4225 18615 4305
rect 18635 4225 18645 4305
rect 18605 4215 18645 4225
rect 18695 4305 18735 4315
rect 18695 4225 18705 4305
rect 18725 4225 18735 4305
rect 18695 4215 18735 4225
rect 18785 4305 18825 4315
rect 18785 4225 18795 4305
rect 18815 4225 18825 4305
rect 18785 4215 18825 4225
rect 18875 4305 18915 4315
rect 18875 4225 18885 4305
rect 18905 4225 18915 4305
rect 18875 4215 18915 4225
rect 18965 4305 19005 4315
rect 18965 4225 18975 4305
rect 18995 4225 19005 4305
rect 18965 4215 19005 4225
rect 19055 4305 19095 4315
rect 19055 4225 19065 4305
rect 19085 4225 19095 4305
rect 19055 4215 19095 4225
rect 19145 4305 19185 4315
rect 19145 4225 19155 4305
rect 19175 4225 19185 4305
rect 19145 4215 19185 4225
rect 19235 4305 19275 4315
rect 19235 4225 19245 4305
rect 19265 4225 19275 4305
rect 19235 4215 19275 4225
rect 19325 4305 19365 4315
rect 19325 4225 19335 4305
rect 19355 4225 19365 4305
rect 19325 4215 19365 4225
rect 19415 4305 19455 4315
rect 19415 4225 19425 4305
rect 19445 4225 19455 4305
rect 19415 4215 19455 4225
rect 19505 4305 19545 4315
rect 19505 4225 19515 4305
rect 19535 4225 19545 4305
rect 19505 4215 19545 4225
rect 19595 4305 19635 4315
rect 19595 4225 19605 4305
rect 19625 4225 19635 4305
rect 19595 4215 19635 4225
rect 19685 4305 19725 4315
rect 19685 4225 19695 4305
rect 19715 4225 19725 4305
rect 19685 4215 19725 4225
rect 19775 4305 19815 4315
rect 19775 4225 19785 4305
rect 19805 4225 19815 4305
rect 19775 4215 19815 4225
rect 19865 4305 19905 4315
rect 19865 4225 19875 4305
rect 19895 4225 19905 4305
rect 19865 4215 19905 4225
rect 19955 4305 19995 4315
rect 19955 4225 19965 4305
rect 19985 4225 19995 4305
rect 19955 4215 19995 4225
rect 20045 4305 20085 4315
rect 20045 4225 20055 4305
rect 20075 4225 20085 4305
rect 20045 4215 20085 4225
rect 20135 4305 20175 4315
rect 20135 4225 20145 4305
rect 20165 4225 20175 4305
rect 20135 4215 20175 4225
rect 20225 4305 20265 4315
rect 20225 4225 20235 4305
rect 20255 4225 20265 4305
rect 20225 4215 20265 4225
rect 20315 4305 20355 4315
rect 20315 4225 20325 4305
rect 20345 4225 20355 4305
rect 20315 4215 20355 4225
rect 20405 4305 20445 4315
rect 20405 4225 20415 4305
rect 20435 4225 20445 4305
rect 20405 4215 20445 4225
rect 20495 4305 20535 4315
rect 20495 4225 20505 4305
rect 20525 4225 20535 4305
rect 20495 4215 20535 4225
rect 20585 4305 20625 4315
rect 20585 4225 20595 4305
rect 20615 4225 20625 4305
rect 20585 4215 20625 4225
rect 20675 4305 20715 4315
rect 20675 4225 20685 4305
rect 20705 4225 20715 4305
rect 20675 4215 20715 4225
<< mvndiffc >>
rect 9165 3485 9185 3565
rect 9255 3485 9275 3565
rect 9345 3485 9365 3565
rect 9435 3485 9455 3565
rect 9525 3485 9545 3565
rect 9615 3485 9635 3565
rect 9705 3485 9725 3565
rect 9795 3485 9815 3565
rect 9885 3485 9905 3565
rect 9975 3485 9995 3565
rect 10065 3485 10085 3565
rect 10155 3485 10175 3565
rect 10245 3485 10265 3565
rect 10335 3485 10355 3565
rect 10425 3485 10445 3565
rect 10515 3485 10535 3565
rect 10605 3485 10625 3565
rect 10695 3485 10715 3565
rect 10785 3485 10805 3565
rect 10875 3485 10895 3565
rect 10965 3485 10985 3565
rect 11055 3485 11075 3565
rect 11145 3485 11165 3565
rect 11235 3485 11255 3565
rect 11325 3485 11345 3565
rect 11415 3485 11435 3565
rect 11505 3485 11525 3565
rect 11595 3485 11615 3565
rect 11685 3485 11705 3565
rect 11775 3485 11795 3565
rect 11865 3485 11885 3565
rect 11955 3485 11975 3565
rect 12045 3485 12065 3565
rect 12135 3485 12155 3565
rect 12225 3485 12245 3565
rect 12315 3485 12335 3565
rect 12405 3485 12425 3565
rect 12495 3485 12515 3565
rect 12585 3485 12605 3565
rect 12675 3485 12695 3565
rect 12765 3485 12785 3565
rect 12855 3485 12875 3565
rect 12945 3485 12965 3565
rect 13035 3485 13055 3565
rect 13125 3485 13145 3565
rect 13215 3485 13235 3565
rect 13305 3485 13325 3565
rect 13395 3485 13415 3565
rect 13485 3485 13505 3565
rect 13575 3485 13595 3565
rect 13665 3485 13685 3565
rect 13755 3485 13775 3565
rect 13845 3485 13865 3565
rect 13935 3485 13955 3565
rect 14025 3485 14045 3565
rect 14115 3485 14135 3565
rect 14205 3485 14225 3565
rect 14295 3485 14315 3565
rect 14385 3485 14405 3565
rect 14475 3485 14495 3565
rect 14565 3485 14585 3565
rect 14655 3485 14675 3565
rect 14745 3485 14765 3565
rect 14835 3485 14855 3565
rect 14925 3485 14945 3565
rect 15015 3485 15035 3565
rect 15105 3485 15125 3565
rect 15195 3485 15215 3565
rect 15285 3485 15305 3565
rect 15375 3485 15395 3565
rect 15465 3485 15485 3565
rect 15555 3485 15575 3565
rect 15645 3485 15665 3565
rect 15735 3485 15755 3565
rect 15825 3485 15845 3565
rect 15915 3485 15935 3565
rect 16005 3485 16025 3565
rect 16095 3485 16115 3565
rect 16185 3485 16205 3565
rect 16275 3485 16295 3565
rect 16365 3485 16385 3565
rect 16455 3485 16475 3565
rect 16545 3485 16565 3565
rect 16635 3485 16655 3565
rect 16725 3485 16745 3565
rect 16815 3485 16835 3565
rect 16905 3485 16925 3565
rect 16995 3485 17015 3565
rect 17085 3485 17105 3565
rect 17175 3485 17195 3565
rect 17265 3485 17285 3565
rect 17355 3485 17375 3565
rect 17445 3485 17465 3565
rect 17535 3485 17555 3565
rect 17625 3485 17645 3565
rect 17715 3485 17735 3565
rect 17805 3485 17825 3565
rect 17895 3485 17915 3565
rect 17985 3485 18005 3565
rect 18075 3485 18095 3565
rect 18165 3485 18185 3565
rect 18255 3485 18275 3565
rect 18345 3485 18365 3565
rect 18435 3485 18455 3565
rect 18525 3485 18545 3565
rect 18615 3485 18635 3565
rect 18705 3485 18725 3565
rect 18795 3485 18815 3565
rect 18885 3485 18905 3565
rect 18975 3485 18995 3565
rect 19065 3485 19085 3565
rect 19155 3485 19175 3565
rect 19245 3485 19265 3565
rect 19335 3485 19355 3565
rect 19425 3485 19445 3565
rect 19515 3485 19535 3565
rect 19605 3485 19625 3565
rect 19695 3485 19715 3565
rect 19785 3485 19805 3565
rect 19875 3485 19895 3565
rect 19965 3485 19985 3565
rect 20055 3485 20075 3565
rect 20145 3485 20165 3565
rect 20235 3485 20255 3565
rect 20325 3485 20345 3565
rect 20415 3485 20435 3565
rect 20505 3485 20525 3565
rect 20595 3485 20615 3565
rect 20685 3485 20705 3565
<< mvpdiffc >>
rect 9165 4225 9185 4305
rect 9255 4225 9275 4305
rect 9345 4225 9365 4305
rect 9435 4225 9455 4305
rect 9525 4225 9545 4305
rect 9615 4225 9635 4305
rect 9705 4225 9725 4305
rect 9795 4225 9815 4305
rect 9885 4225 9905 4305
rect 9975 4225 9995 4305
rect 10065 4225 10085 4305
rect 10155 4225 10175 4305
rect 10245 4225 10265 4305
rect 10335 4225 10355 4305
rect 10425 4225 10445 4305
rect 10515 4225 10535 4305
rect 10605 4225 10625 4305
rect 10695 4225 10715 4305
rect 10785 4225 10805 4305
rect 10875 4225 10895 4305
rect 10965 4225 10985 4305
rect 11055 4225 11075 4305
rect 11145 4225 11165 4305
rect 11235 4225 11255 4305
rect 11325 4225 11345 4305
rect 11415 4225 11435 4305
rect 11505 4225 11525 4305
rect 11595 4225 11615 4305
rect 11685 4225 11705 4305
rect 11775 4225 11795 4305
rect 11865 4225 11885 4305
rect 11955 4225 11975 4305
rect 12045 4225 12065 4305
rect 12135 4225 12155 4305
rect 12225 4225 12245 4305
rect 12315 4225 12335 4305
rect 12405 4225 12425 4305
rect 12495 4225 12515 4305
rect 12585 4225 12605 4305
rect 12675 4225 12695 4305
rect 12765 4225 12785 4305
rect 12855 4225 12875 4305
rect 12945 4225 12965 4305
rect 13035 4225 13055 4305
rect 13125 4225 13145 4305
rect 13215 4225 13235 4305
rect 13305 4225 13325 4305
rect 13395 4225 13415 4305
rect 13485 4225 13505 4305
rect 13575 4225 13595 4305
rect 13665 4225 13685 4305
rect 13755 4225 13775 4305
rect 13845 4225 13865 4305
rect 13935 4225 13955 4305
rect 14025 4225 14045 4305
rect 14115 4225 14135 4305
rect 14205 4225 14225 4305
rect 14295 4225 14315 4305
rect 14385 4225 14405 4305
rect 14475 4225 14495 4305
rect 14565 4225 14585 4305
rect 14655 4225 14675 4305
rect 14745 4225 14765 4305
rect 14835 4225 14855 4305
rect 14925 4225 14945 4305
rect 15015 4225 15035 4305
rect 15105 4225 15125 4305
rect 15195 4225 15215 4305
rect 15285 4225 15305 4305
rect 15375 4225 15395 4305
rect 15465 4225 15485 4305
rect 15555 4225 15575 4305
rect 15645 4225 15665 4305
rect 15735 4225 15755 4305
rect 15825 4225 15845 4305
rect 15915 4225 15935 4305
rect 16005 4225 16025 4305
rect 16095 4225 16115 4305
rect 16185 4225 16205 4305
rect 16275 4225 16295 4305
rect 16365 4225 16385 4305
rect 16455 4225 16475 4305
rect 16545 4225 16565 4305
rect 16635 4225 16655 4305
rect 16725 4225 16745 4305
rect 16815 4225 16835 4305
rect 16905 4225 16925 4305
rect 16995 4225 17015 4305
rect 17085 4225 17105 4305
rect 17175 4225 17195 4305
rect 17265 4225 17285 4305
rect 17355 4225 17375 4305
rect 17445 4225 17465 4305
rect 17535 4225 17555 4305
rect 17625 4225 17645 4305
rect 17715 4225 17735 4305
rect 17805 4225 17825 4305
rect 17895 4225 17915 4305
rect 17985 4225 18005 4305
rect 18075 4225 18095 4305
rect 18165 4225 18185 4305
rect 18255 4225 18275 4305
rect 18345 4225 18365 4305
rect 18435 4225 18455 4305
rect 18525 4225 18545 4305
rect 18615 4225 18635 4305
rect 18705 4225 18725 4305
rect 18795 4225 18815 4305
rect 18885 4225 18905 4305
rect 18975 4225 18995 4305
rect 19065 4225 19085 4305
rect 19155 4225 19175 4305
rect 19245 4225 19265 4305
rect 19335 4225 19355 4305
rect 19425 4225 19445 4305
rect 19515 4225 19535 4305
rect 19605 4225 19625 4305
rect 19695 4225 19715 4305
rect 19785 4225 19805 4305
rect 19875 4225 19895 4305
rect 19965 4225 19985 4305
rect 20055 4225 20075 4305
rect 20145 4225 20165 4305
rect 20235 4225 20255 4305
rect 20325 4225 20345 4305
rect 20415 4225 20435 4305
rect 20505 4225 20525 4305
rect 20595 4225 20615 4305
rect 20685 4225 20705 4305
<< psubdiff >>
rect 9030 4065 9050 4375
rect 20820 4065 20840 4375
rect 9030 4045 9210 4065
rect 9230 4045 9300 4065
rect 9320 4045 9390 4065
rect 9410 4045 9480 4065
rect 9500 4045 9570 4065
rect 9590 4045 9660 4065
rect 9680 4045 9750 4065
rect 9770 4045 9840 4065
rect 9860 4045 9930 4065
rect 9950 4045 10020 4065
rect 10040 4045 10110 4065
rect 10130 4045 10200 4065
rect 10220 4045 10290 4065
rect 10310 4045 10380 4065
rect 10400 4045 10470 4065
rect 10490 4045 10560 4065
rect 10580 4045 10650 4065
rect 10670 4045 10740 4065
rect 10760 4045 10830 4065
rect 10850 4045 10920 4065
rect 10940 4045 11010 4065
rect 11030 4045 11100 4065
rect 11120 4045 11190 4065
rect 11210 4045 11280 4065
rect 11300 4045 11370 4065
rect 11390 4045 11460 4065
rect 11480 4045 11550 4065
rect 11570 4045 11640 4065
rect 11660 4045 11730 4065
rect 11750 4045 11820 4065
rect 11840 4045 11910 4065
rect 11930 4045 12000 4065
rect 12020 4045 12090 4065
rect 12110 4045 12180 4065
rect 12200 4045 12270 4065
rect 12290 4045 12360 4065
rect 12380 4045 12450 4065
rect 12470 4045 12540 4065
rect 12560 4045 12630 4065
rect 12650 4045 12720 4065
rect 12740 4045 12810 4065
rect 12830 4045 12900 4065
rect 12920 4045 12990 4065
rect 13010 4045 13080 4065
rect 13100 4045 13170 4065
rect 13190 4045 13260 4065
rect 13280 4045 13350 4065
rect 13370 4045 13440 4065
rect 13460 4045 13530 4065
rect 13550 4045 13620 4065
rect 13640 4045 13710 4065
rect 13730 4045 13800 4065
rect 13820 4045 13890 4065
rect 13910 4045 13980 4065
rect 14000 4045 14070 4065
rect 14090 4045 14160 4065
rect 14180 4045 14250 4065
rect 14270 4045 14340 4065
rect 14360 4045 14430 4065
rect 14450 4045 14520 4065
rect 14540 4045 14610 4065
rect 14630 4045 14700 4065
rect 14720 4045 14790 4065
rect 14810 4045 14880 4065
rect 14900 4045 14970 4065
rect 14990 4045 15060 4065
rect 15080 4045 15150 4065
rect 15170 4045 15240 4065
rect 15260 4045 15330 4065
rect 15350 4045 15420 4065
rect 15440 4045 15510 4065
rect 15530 4045 15600 4065
rect 15620 4045 15690 4065
rect 15710 4045 15780 4065
rect 15800 4045 15870 4065
rect 15890 4045 15960 4065
rect 15980 4045 16050 4065
rect 16070 4045 16140 4065
rect 16160 4045 16230 4065
rect 16250 4045 16320 4065
rect 16340 4045 16410 4065
rect 16430 4045 16500 4065
rect 16520 4045 16590 4065
rect 16610 4045 16680 4065
rect 16700 4045 16770 4065
rect 16790 4045 16860 4065
rect 16880 4045 16950 4065
rect 16970 4045 17040 4065
rect 17060 4045 17130 4065
rect 17150 4045 17220 4065
rect 17240 4045 17310 4065
rect 17330 4045 17400 4065
rect 17420 4045 17490 4065
rect 17510 4045 17580 4065
rect 17600 4045 17670 4065
rect 17690 4045 17760 4065
rect 17780 4045 17850 4065
rect 17870 4045 17940 4065
rect 17960 4045 18030 4065
rect 18050 4045 18120 4065
rect 18140 4045 18210 4065
rect 18230 4045 18300 4065
rect 18320 4045 18390 4065
rect 18410 4045 18480 4065
rect 18500 4045 18570 4065
rect 18590 4045 18660 4065
rect 18680 4045 18750 4065
rect 18770 4045 18840 4065
rect 18860 4045 18930 4065
rect 18950 4045 19020 4065
rect 19040 4045 19110 4065
rect 19130 4045 19200 4065
rect 19220 4045 19290 4065
rect 19310 4045 19380 4065
rect 19400 4045 19470 4065
rect 19490 4045 19560 4065
rect 19580 4045 19650 4065
rect 19670 4045 19740 4065
rect 19760 4045 19830 4065
rect 19850 4045 19920 4065
rect 19940 4045 20010 4065
rect 20030 4045 20100 4065
rect 20120 4045 20190 4065
rect 20210 4045 20280 4065
rect 20300 4045 20370 4065
rect 20390 4045 20460 4065
rect 20480 4045 20550 4065
rect 20570 4045 20640 4065
rect 20660 4045 20840 4065
rect 9030 3645 9210 3665
rect 9230 3645 9300 3665
rect 9320 3645 9390 3665
rect 9410 3645 9480 3665
rect 9500 3645 9570 3665
rect 9590 3645 9660 3665
rect 9680 3645 9750 3665
rect 9770 3645 9840 3665
rect 9860 3645 9930 3665
rect 9950 3645 10020 3665
rect 10040 3645 10110 3665
rect 10130 3645 10200 3665
rect 10220 3645 10290 3665
rect 10310 3645 10380 3665
rect 10400 3645 10470 3665
rect 10490 3645 10560 3665
rect 10580 3645 10650 3665
rect 10670 3645 10740 3665
rect 10760 3645 10830 3665
rect 10850 3645 10920 3665
rect 10940 3645 11010 3665
rect 11030 3645 11100 3665
rect 11120 3645 11190 3665
rect 11210 3645 11280 3665
rect 11300 3645 11370 3665
rect 11390 3645 11460 3665
rect 11480 3645 11550 3665
rect 11570 3645 11640 3665
rect 11660 3645 11730 3665
rect 11750 3645 11820 3665
rect 11840 3645 11910 3665
rect 11930 3645 12000 3665
rect 12020 3645 12090 3665
rect 12110 3645 12180 3665
rect 12200 3645 12270 3665
rect 12290 3645 12360 3665
rect 12380 3645 12450 3665
rect 12470 3645 12540 3665
rect 12560 3645 12630 3665
rect 12650 3645 12720 3665
rect 12740 3645 12810 3665
rect 12830 3645 12900 3665
rect 12920 3645 12990 3665
rect 13010 3645 13080 3665
rect 13100 3645 13170 3665
rect 13190 3645 13260 3665
rect 13280 3645 13350 3665
rect 13370 3645 13440 3665
rect 13460 3645 13530 3665
rect 13550 3645 13620 3665
rect 13640 3645 13710 3665
rect 13730 3645 13800 3665
rect 13820 3645 13890 3665
rect 13910 3645 13980 3665
rect 14000 3645 14070 3665
rect 14090 3645 14160 3665
rect 14180 3645 14250 3665
rect 14270 3645 14340 3665
rect 14360 3645 14430 3665
rect 14450 3645 14520 3665
rect 14540 3645 14610 3665
rect 14630 3645 14700 3665
rect 14720 3645 14790 3665
rect 14810 3645 14880 3665
rect 14900 3645 14970 3665
rect 14990 3645 15060 3665
rect 15080 3645 15150 3665
rect 15170 3645 15240 3665
rect 15260 3645 15330 3665
rect 15350 3645 15420 3665
rect 15440 3645 15510 3665
rect 15530 3645 15600 3665
rect 15620 3645 15690 3665
rect 15710 3645 15780 3665
rect 15800 3645 15870 3665
rect 15890 3645 15960 3665
rect 15980 3645 16050 3665
rect 16070 3645 16140 3665
rect 16160 3645 16230 3665
rect 16250 3645 16320 3665
rect 16340 3645 16410 3665
rect 16430 3645 16500 3665
rect 16520 3645 16590 3665
rect 16610 3645 16680 3665
rect 16700 3645 16770 3665
rect 16790 3645 16860 3665
rect 16880 3645 16950 3665
rect 16970 3645 17040 3665
rect 17060 3645 17130 3665
rect 17150 3645 17220 3665
rect 17240 3645 17310 3665
rect 17330 3645 17400 3665
rect 17420 3645 17490 3665
rect 17510 3645 17580 3665
rect 17600 3645 17670 3665
rect 17690 3645 17760 3665
rect 17780 3645 17850 3665
rect 17870 3645 17940 3665
rect 17960 3645 18030 3665
rect 18050 3645 18120 3665
rect 18140 3645 18210 3665
rect 18230 3645 18300 3665
rect 18320 3645 18390 3665
rect 18410 3645 18480 3665
rect 18500 3645 18570 3665
rect 18590 3645 18660 3665
rect 18680 3645 18750 3665
rect 18770 3645 18840 3665
rect 18860 3645 18930 3665
rect 18950 3645 19020 3665
rect 19040 3645 19110 3665
rect 19130 3645 19200 3665
rect 19220 3645 19290 3665
rect 19310 3645 19380 3665
rect 19400 3645 19470 3665
rect 19490 3645 19560 3665
rect 19580 3645 19650 3665
rect 19670 3645 19740 3665
rect 19760 3645 19830 3665
rect 19850 3645 19920 3665
rect 19940 3645 20010 3665
rect 20030 3645 20100 3665
rect 20120 3645 20190 3665
rect 20210 3645 20280 3665
rect 20300 3645 20370 3665
rect 20390 3645 20460 3665
rect 20480 3645 20550 3665
rect 20570 3645 20640 3665
rect 20660 3645 20840 3665
rect 9030 3445 9050 3645
rect 20820 3445 20840 3645
rect 9020 3425 9210 3445
rect 9230 3425 9300 3445
rect 9320 3425 9390 3445
rect 9410 3425 9480 3445
rect 9500 3425 9570 3445
rect 9590 3425 9660 3445
rect 9680 3425 9750 3445
rect 9770 3425 9840 3445
rect 9860 3425 9930 3445
rect 9950 3425 10020 3445
rect 10040 3425 10110 3445
rect 10130 3425 10200 3445
rect 10220 3425 10290 3445
rect 10310 3425 10380 3445
rect 10400 3425 10470 3445
rect 10490 3425 10560 3445
rect 10580 3425 10650 3445
rect 10670 3425 10740 3445
rect 10760 3425 10830 3445
rect 10850 3425 10920 3445
rect 10940 3425 11010 3445
rect 11030 3425 11100 3445
rect 11120 3425 11190 3445
rect 11210 3425 11280 3445
rect 11300 3425 11370 3445
rect 11390 3425 11460 3445
rect 11480 3425 11550 3445
rect 11570 3425 11640 3445
rect 11660 3425 11730 3445
rect 11750 3425 11820 3445
rect 11840 3425 11910 3445
rect 11930 3425 12000 3445
rect 12020 3425 12090 3445
rect 12110 3425 12180 3445
rect 12200 3425 12270 3445
rect 12290 3425 12360 3445
rect 12380 3425 12450 3445
rect 12470 3425 12540 3445
rect 12560 3425 12630 3445
rect 12650 3425 12720 3445
rect 12740 3425 12810 3445
rect 12830 3425 12900 3445
rect 12920 3425 12990 3445
rect 13010 3425 13080 3445
rect 13100 3425 13170 3445
rect 13190 3425 13260 3445
rect 13280 3425 13350 3445
rect 13370 3425 13440 3445
rect 13460 3425 13530 3445
rect 13550 3425 13620 3445
rect 13640 3425 13710 3445
rect 13730 3425 13800 3445
rect 13820 3425 13890 3445
rect 13910 3425 13980 3445
rect 14000 3425 14070 3445
rect 14090 3425 14160 3445
rect 14180 3425 14250 3445
rect 14270 3425 14340 3445
rect 14360 3425 14430 3445
rect 14450 3425 14520 3445
rect 14540 3425 14610 3445
rect 14630 3425 14700 3445
rect 14720 3425 14790 3445
rect 14810 3425 14880 3445
rect 14900 3425 14970 3445
rect 14990 3425 15060 3445
rect 15080 3425 15150 3445
rect 15170 3425 15240 3445
rect 15260 3425 15330 3445
rect 15350 3425 15420 3445
rect 15440 3425 15510 3445
rect 15530 3425 15600 3445
rect 15620 3425 15690 3445
rect 15710 3425 15780 3445
rect 15800 3425 15870 3445
rect 15890 3425 15960 3445
rect 15980 3425 16050 3445
rect 16070 3425 16140 3445
rect 16160 3425 16230 3445
rect 16250 3425 16320 3445
rect 16340 3425 16410 3445
rect 16430 3425 16500 3445
rect 16520 3425 16590 3445
rect 16610 3425 16680 3445
rect 16700 3425 16770 3445
rect 16790 3425 16860 3445
rect 16880 3425 16950 3445
rect 16970 3425 17040 3445
rect 17060 3425 17130 3445
rect 17150 3425 17220 3445
rect 17240 3425 17310 3445
rect 17330 3425 17400 3445
rect 17420 3425 17490 3445
rect 17510 3425 17580 3445
rect 17600 3425 17670 3445
rect 17690 3425 17760 3445
rect 17780 3425 17850 3445
rect 17870 3425 17940 3445
rect 17960 3425 18030 3445
rect 18050 3425 18120 3445
rect 18140 3425 18210 3445
rect 18230 3425 18300 3445
rect 18320 3425 18390 3445
rect 18410 3425 18480 3445
rect 18500 3425 18570 3445
rect 18590 3425 18660 3445
rect 18680 3425 18750 3445
rect 18770 3425 18840 3445
rect 18860 3425 18930 3445
rect 18950 3425 19020 3445
rect 19040 3425 19110 3445
rect 19130 3425 19200 3445
rect 19220 3425 19290 3445
rect 19310 3425 19380 3445
rect 19400 3425 19470 3445
rect 19490 3425 19560 3445
rect 19580 3425 19650 3445
rect 19670 3425 19740 3445
rect 19760 3425 19830 3445
rect 19850 3425 19920 3445
rect 19940 3425 20010 3445
rect 20030 3425 20100 3445
rect 20120 3425 20190 3445
rect 20210 3425 20280 3445
rect 20300 3425 20370 3445
rect 20390 3425 20460 3445
rect 20480 3425 20550 3445
rect 20570 3425 20640 3445
rect 20660 3425 20850 3445
<< nsubdiff >>
rect 9105 4345 9210 4365
rect 9230 4345 9300 4365
rect 9320 4345 9390 4365
rect 9410 4345 9480 4365
rect 9500 4345 9570 4365
rect 9590 4345 9660 4365
rect 9680 4345 9750 4365
rect 9770 4345 9840 4365
rect 9860 4345 9930 4365
rect 9950 4345 10020 4365
rect 10040 4345 10110 4365
rect 10130 4345 10200 4365
rect 10220 4345 10290 4365
rect 10310 4345 10380 4365
rect 10400 4345 10470 4365
rect 10490 4345 10560 4365
rect 10580 4345 10650 4365
rect 10670 4345 10740 4365
rect 10760 4345 10830 4365
rect 10850 4345 10920 4365
rect 10940 4345 11010 4365
rect 11030 4345 11100 4365
rect 11120 4345 11190 4365
rect 11210 4345 11280 4365
rect 11300 4345 11370 4365
rect 11390 4345 11460 4365
rect 11480 4345 11550 4365
rect 11570 4345 11640 4365
rect 11660 4345 11730 4365
rect 11750 4345 11820 4365
rect 11840 4345 11910 4365
rect 11930 4345 12000 4365
rect 12020 4345 12090 4365
rect 12110 4345 12180 4365
rect 12200 4345 12270 4365
rect 12290 4345 12360 4365
rect 12380 4345 12450 4365
rect 12470 4345 12540 4365
rect 12560 4345 12630 4365
rect 12650 4345 12720 4365
rect 12740 4345 12810 4365
rect 12830 4345 12900 4365
rect 12920 4345 12990 4365
rect 13010 4345 13080 4365
rect 13100 4345 13170 4365
rect 13190 4345 13260 4365
rect 13280 4345 13350 4365
rect 13370 4345 13440 4365
rect 13460 4345 13530 4365
rect 13550 4345 13620 4365
rect 13640 4345 13710 4365
rect 13730 4345 13800 4365
rect 13820 4345 13890 4365
rect 13910 4345 13980 4365
rect 14000 4345 14070 4365
rect 14090 4345 14160 4365
rect 14180 4345 14250 4365
rect 14270 4345 14340 4365
rect 14360 4345 14430 4365
rect 14450 4345 14520 4365
rect 14540 4345 14610 4365
rect 14630 4345 14700 4365
rect 14720 4345 14790 4365
rect 14810 4345 14880 4365
rect 14900 4345 14970 4365
rect 14990 4345 15060 4365
rect 15080 4345 15150 4365
rect 15170 4345 15240 4365
rect 15260 4345 15330 4365
rect 15350 4345 15420 4365
rect 15440 4345 15510 4365
rect 15530 4345 15600 4365
rect 15620 4345 15690 4365
rect 15710 4345 15780 4365
rect 15800 4345 15870 4365
rect 15890 4345 15960 4365
rect 15980 4345 16050 4365
rect 16070 4345 16140 4365
rect 16160 4345 16230 4365
rect 16250 4345 16320 4365
rect 16340 4345 16410 4365
rect 16430 4345 16500 4365
rect 16520 4345 16590 4365
rect 16610 4345 16680 4365
rect 16700 4345 16770 4365
rect 16790 4345 16860 4365
rect 16880 4345 16950 4365
rect 16970 4345 17040 4365
rect 17060 4345 17130 4365
rect 17150 4345 17220 4365
rect 17240 4345 17310 4365
rect 17330 4345 17400 4365
rect 17420 4345 17490 4365
rect 17510 4345 17580 4365
rect 17600 4345 17670 4365
rect 17690 4345 17760 4365
rect 17780 4345 17850 4365
rect 17870 4345 17940 4365
rect 17960 4345 18030 4365
rect 18050 4345 18120 4365
rect 18140 4345 18210 4365
rect 18230 4345 18300 4365
rect 18320 4345 18390 4365
rect 18410 4345 18480 4365
rect 18500 4345 18570 4365
rect 18590 4345 18660 4365
rect 18680 4345 18750 4365
rect 18770 4345 18840 4365
rect 18860 4345 18930 4365
rect 18950 4345 19020 4365
rect 19040 4345 19110 4365
rect 19130 4345 19200 4365
rect 19220 4345 19290 4365
rect 19310 4345 19380 4365
rect 19400 4345 19470 4365
rect 19490 4345 19560 4365
rect 19580 4345 19650 4365
rect 19670 4345 19740 4365
rect 19760 4345 19830 4365
rect 19850 4345 19920 4365
rect 19940 4345 20010 4365
rect 20030 4345 20100 4365
rect 20120 4345 20190 4365
rect 20210 4345 20280 4365
rect 20300 4345 20370 4365
rect 20390 4345 20460 4365
rect 20480 4345 20550 4365
rect 20570 4345 20640 4365
rect 20660 4345 20765 4365
rect 9105 4145 9125 4345
rect 20745 4145 20765 4345
rect 9105 4125 9210 4145
rect 9230 4125 9300 4145
rect 9320 4125 9390 4145
rect 9410 4125 9480 4145
rect 9500 4125 9570 4145
rect 9590 4125 9660 4145
rect 9680 4125 9750 4145
rect 9770 4125 9840 4145
rect 9860 4125 9930 4145
rect 9950 4125 10020 4145
rect 10040 4125 10110 4145
rect 10130 4125 10200 4145
rect 10220 4125 10290 4145
rect 10310 4125 10380 4145
rect 10400 4125 10470 4145
rect 10490 4125 10560 4145
rect 10580 4125 10650 4145
rect 10670 4125 10740 4145
rect 10760 4125 10830 4145
rect 10850 4125 10920 4145
rect 10940 4125 11010 4145
rect 11030 4125 11100 4145
rect 11120 4125 11190 4145
rect 11210 4125 11280 4145
rect 11300 4125 11370 4145
rect 11390 4125 11460 4145
rect 11480 4125 11550 4145
rect 11570 4125 11640 4145
rect 11660 4125 11730 4145
rect 11750 4125 11820 4145
rect 11840 4125 11910 4145
rect 11930 4125 12000 4145
rect 12020 4125 12090 4145
rect 12110 4125 12180 4145
rect 12200 4125 12270 4145
rect 12290 4125 12360 4145
rect 12380 4125 12450 4145
rect 12470 4125 12540 4145
rect 12560 4125 12630 4145
rect 12650 4125 12720 4145
rect 12740 4125 12810 4145
rect 12830 4125 12900 4145
rect 12920 4125 12990 4145
rect 13010 4125 13080 4145
rect 13100 4125 13170 4145
rect 13190 4125 13260 4145
rect 13280 4125 13350 4145
rect 13370 4125 13440 4145
rect 13460 4125 13530 4145
rect 13550 4125 13620 4145
rect 13640 4125 13710 4145
rect 13730 4125 13800 4145
rect 13820 4125 13890 4145
rect 13910 4125 13980 4145
rect 14000 4125 14070 4145
rect 14090 4125 14160 4145
rect 14180 4125 14250 4145
rect 14270 4125 14340 4145
rect 14360 4125 14430 4145
rect 14450 4125 14520 4145
rect 14540 4125 14610 4145
rect 14630 4125 14700 4145
rect 14720 4125 14790 4145
rect 14810 4125 14880 4145
rect 14900 4125 14970 4145
rect 14990 4125 15060 4145
rect 15080 4125 15150 4145
rect 15170 4125 15240 4145
rect 15260 4125 15330 4145
rect 15350 4125 15420 4145
rect 15440 4125 15510 4145
rect 15530 4125 15600 4145
rect 15620 4125 15690 4145
rect 15710 4125 15780 4145
rect 15800 4125 15870 4145
rect 15890 4125 15960 4145
rect 15980 4125 16050 4145
rect 16070 4125 16140 4145
rect 16160 4125 16230 4145
rect 16250 4125 16320 4145
rect 16340 4125 16410 4145
rect 16430 4125 16500 4145
rect 16520 4125 16590 4145
rect 16610 4125 16680 4145
rect 16700 4125 16770 4145
rect 16790 4125 16860 4145
rect 16880 4125 16950 4145
rect 16970 4125 17040 4145
rect 17060 4125 17130 4145
rect 17150 4125 17220 4145
rect 17240 4125 17310 4145
rect 17330 4125 17400 4145
rect 17420 4125 17490 4145
rect 17510 4125 17580 4145
rect 17600 4125 17670 4145
rect 17690 4125 17760 4145
rect 17780 4125 17850 4145
rect 17870 4125 17940 4145
rect 17960 4125 18030 4145
rect 18050 4125 18120 4145
rect 18140 4125 18210 4145
rect 18230 4125 18300 4145
rect 18320 4125 18390 4145
rect 18410 4125 18480 4145
rect 18500 4125 18570 4145
rect 18590 4125 18660 4145
rect 18680 4125 18750 4145
rect 18770 4125 18840 4145
rect 18860 4125 18930 4145
rect 18950 4125 19020 4145
rect 19040 4125 19110 4145
rect 19130 4125 19200 4145
rect 19220 4125 19290 4145
rect 19310 4125 19380 4145
rect 19400 4125 19470 4145
rect 19490 4125 19560 4145
rect 19580 4125 19650 4145
rect 19670 4125 19740 4145
rect 19760 4125 19830 4145
rect 19850 4125 19920 4145
rect 19940 4125 20010 4145
rect 20030 4125 20100 4145
rect 20120 4125 20190 4145
rect 20210 4125 20280 4145
rect 20300 4125 20370 4145
rect 20390 4125 20460 4145
rect 20480 4125 20550 4145
rect 20570 4125 20640 4145
rect 20660 4125 20765 4145
<< psubdiffcont >>
rect 9210 4045 9230 4065
rect 9300 4045 9320 4065
rect 9390 4045 9410 4065
rect 9480 4045 9500 4065
rect 9570 4045 9590 4065
rect 9660 4045 9680 4065
rect 9750 4045 9770 4065
rect 9840 4045 9860 4065
rect 9930 4045 9950 4065
rect 10020 4045 10040 4065
rect 10110 4045 10130 4065
rect 10200 4045 10220 4065
rect 10290 4045 10310 4065
rect 10380 4045 10400 4065
rect 10470 4045 10490 4065
rect 10560 4045 10580 4065
rect 10650 4045 10670 4065
rect 10740 4045 10760 4065
rect 10830 4045 10850 4065
rect 10920 4045 10940 4065
rect 11010 4045 11030 4065
rect 11100 4045 11120 4065
rect 11190 4045 11210 4065
rect 11280 4045 11300 4065
rect 11370 4045 11390 4065
rect 11460 4045 11480 4065
rect 11550 4045 11570 4065
rect 11640 4045 11660 4065
rect 11730 4045 11750 4065
rect 11820 4045 11840 4065
rect 11910 4045 11930 4065
rect 12000 4045 12020 4065
rect 12090 4045 12110 4065
rect 12180 4045 12200 4065
rect 12270 4045 12290 4065
rect 12360 4045 12380 4065
rect 12450 4045 12470 4065
rect 12540 4045 12560 4065
rect 12630 4045 12650 4065
rect 12720 4045 12740 4065
rect 12810 4045 12830 4065
rect 12900 4045 12920 4065
rect 12990 4045 13010 4065
rect 13080 4045 13100 4065
rect 13170 4045 13190 4065
rect 13260 4045 13280 4065
rect 13350 4045 13370 4065
rect 13440 4045 13460 4065
rect 13530 4045 13550 4065
rect 13620 4045 13640 4065
rect 13710 4045 13730 4065
rect 13800 4045 13820 4065
rect 13890 4045 13910 4065
rect 13980 4045 14000 4065
rect 14070 4045 14090 4065
rect 14160 4045 14180 4065
rect 14250 4045 14270 4065
rect 14340 4045 14360 4065
rect 14430 4045 14450 4065
rect 14520 4045 14540 4065
rect 14610 4045 14630 4065
rect 14700 4045 14720 4065
rect 14790 4045 14810 4065
rect 14880 4045 14900 4065
rect 14970 4045 14990 4065
rect 15060 4045 15080 4065
rect 15150 4045 15170 4065
rect 15240 4045 15260 4065
rect 15330 4045 15350 4065
rect 15420 4045 15440 4065
rect 15510 4045 15530 4065
rect 15600 4045 15620 4065
rect 15690 4045 15710 4065
rect 15780 4045 15800 4065
rect 15870 4045 15890 4065
rect 15960 4045 15980 4065
rect 16050 4045 16070 4065
rect 16140 4045 16160 4065
rect 16230 4045 16250 4065
rect 16320 4045 16340 4065
rect 16410 4045 16430 4065
rect 16500 4045 16520 4065
rect 16590 4045 16610 4065
rect 16680 4045 16700 4065
rect 16770 4045 16790 4065
rect 16860 4045 16880 4065
rect 16950 4045 16970 4065
rect 17040 4045 17060 4065
rect 17130 4045 17150 4065
rect 17220 4045 17240 4065
rect 17310 4045 17330 4065
rect 17400 4045 17420 4065
rect 17490 4045 17510 4065
rect 17580 4045 17600 4065
rect 17670 4045 17690 4065
rect 17760 4045 17780 4065
rect 17850 4045 17870 4065
rect 17940 4045 17960 4065
rect 18030 4045 18050 4065
rect 18120 4045 18140 4065
rect 18210 4045 18230 4065
rect 18300 4045 18320 4065
rect 18390 4045 18410 4065
rect 18480 4045 18500 4065
rect 18570 4045 18590 4065
rect 18660 4045 18680 4065
rect 18750 4045 18770 4065
rect 18840 4045 18860 4065
rect 18930 4045 18950 4065
rect 19020 4045 19040 4065
rect 19110 4045 19130 4065
rect 19200 4045 19220 4065
rect 19290 4045 19310 4065
rect 19380 4045 19400 4065
rect 19470 4045 19490 4065
rect 19560 4045 19580 4065
rect 19650 4045 19670 4065
rect 19740 4045 19760 4065
rect 19830 4045 19850 4065
rect 19920 4045 19940 4065
rect 20010 4045 20030 4065
rect 20100 4045 20120 4065
rect 20190 4045 20210 4065
rect 20280 4045 20300 4065
rect 20370 4045 20390 4065
rect 20460 4045 20480 4065
rect 20550 4045 20570 4065
rect 20640 4045 20660 4065
rect 9210 3645 9230 3665
rect 9300 3645 9320 3665
rect 9390 3645 9410 3665
rect 9480 3645 9500 3665
rect 9570 3645 9590 3665
rect 9660 3645 9680 3665
rect 9750 3645 9770 3665
rect 9840 3645 9860 3665
rect 9930 3645 9950 3665
rect 10020 3645 10040 3665
rect 10110 3645 10130 3665
rect 10200 3645 10220 3665
rect 10290 3645 10310 3665
rect 10380 3645 10400 3665
rect 10470 3645 10490 3665
rect 10560 3645 10580 3665
rect 10650 3645 10670 3665
rect 10740 3645 10760 3665
rect 10830 3645 10850 3665
rect 10920 3645 10940 3665
rect 11010 3645 11030 3665
rect 11100 3645 11120 3665
rect 11190 3645 11210 3665
rect 11280 3645 11300 3665
rect 11370 3645 11390 3665
rect 11460 3645 11480 3665
rect 11550 3645 11570 3665
rect 11640 3645 11660 3665
rect 11730 3645 11750 3665
rect 11820 3645 11840 3665
rect 11910 3645 11930 3665
rect 12000 3645 12020 3665
rect 12090 3645 12110 3665
rect 12180 3645 12200 3665
rect 12270 3645 12290 3665
rect 12360 3645 12380 3665
rect 12450 3645 12470 3665
rect 12540 3645 12560 3665
rect 12630 3645 12650 3665
rect 12720 3645 12740 3665
rect 12810 3645 12830 3665
rect 12900 3645 12920 3665
rect 12990 3645 13010 3665
rect 13080 3645 13100 3665
rect 13170 3645 13190 3665
rect 13260 3645 13280 3665
rect 13350 3645 13370 3665
rect 13440 3645 13460 3665
rect 13530 3645 13550 3665
rect 13620 3645 13640 3665
rect 13710 3645 13730 3665
rect 13800 3645 13820 3665
rect 13890 3645 13910 3665
rect 13980 3645 14000 3665
rect 14070 3645 14090 3665
rect 14160 3645 14180 3665
rect 14250 3645 14270 3665
rect 14340 3645 14360 3665
rect 14430 3645 14450 3665
rect 14520 3645 14540 3665
rect 14610 3645 14630 3665
rect 14700 3645 14720 3665
rect 14790 3645 14810 3665
rect 14880 3645 14900 3665
rect 14970 3645 14990 3665
rect 15060 3645 15080 3665
rect 15150 3645 15170 3665
rect 15240 3645 15260 3665
rect 15330 3645 15350 3665
rect 15420 3645 15440 3665
rect 15510 3645 15530 3665
rect 15600 3645 15620 3665
rect 15690 3645 15710 3665
rect 15780 3645 15800 3665
rect 15870 3645 15890 3665
rect 15960 3645 15980 3665
rect 16050 3645 16070 3665
rect 16140 3645 16160 3665
rect 16230 3645 16250 3665
rect 16320 3645 16340 3665
rect 16410 3645 16430 3665
rect 16500 3645 16520 3665
rect 16590 3645 16610 3665
rect 16680 3645 16700 3665
rect 16770 3645 16790 3665
rect 16860 3645 16880 3665
rect 16950 3645 16970 3665
rect 17040 3645 17060 3665
rect 17130 3645 17150 3665
rect 17220 3645 17240 3665
rect 17310 3645 17330 3665
rect 17400 3645 17420 3665
rect 17490 3645 17510 3665
rect 17580 3645 17600 3665
rect 17670 3645 17690 3665
rect 17760 3645 17780 3665
rect 17850 3645 17870 3665
rect 17940 3645 17960 3665
rect 18030 3645 18050 3665
rect 18120 3645 18140 3665
rect 18210 3645 18230 3665
rect 18300 3645 18320 3665
rect 18390 3645 18410 3665
rect 18480 3645 18500 3665
rect 18570 3645 18590 3665
rect 18660 3645 18680 3665
rect 18750 3645 18770 3665
rect 18840 3645 18860 3665
rect 18930 3645 18950 3665
rect 19020 3645 19040 3665
rect 19110 3645 19130 3665
rect 19200 3645 19220 3665
rect 19290 3645 19310 3665
rect 19380 3645 19400 3665
rect 19470 3645 19490 3665
rect 19560 3645 19580 3665
rect 19650 3645 19670 3665
rect 19740 3645 19760 3665
rect 19830 3645 19850 3665
rect 19920 3645 19940 3665
rect 20010 3645 20030 3665
rect 20100 3645 20120 3665
rect 20190 3645 20210 3665
rect 20280 3645 20300 3665
rect 20370 3645 20390 3665
rect 20460 3645 20480 3665
rect 20550 3645 20570 3665
rect 20640 3645 20660 3665
rect 9210 3425 9230 3445
rect 9300 3425 9320 3445
rect 9390 3425 9410 3445
rect 9480 3425 9500 3445
rect 9570 3425 9590 3445
rect 9660 3425 9680 3445
rect 9750 3425 9770 3445
rect 9840 3425 9860 3445
rect 9930 3425 9950 3445
rect 10020 3425 10040 3445
rect 10110 3425 10130 3445
rect 10200 3425 10220 3445
rect 10290 3425 10310 3445
rect 10380 3425 10400 3445
rect 10470 3425 10490 3445
rect 10560 3425 10580 3445
rect 10650 3425 10670 3445
rect 10740 3425 10760 3445
rect 10830 3425 10850 3445
rect 10920 3425 10940 3445
rect 11010 3425 11030 3445
rect 11100 3425 11120 3445
rect 11190 3425 11210 3445
rect 11280 3425 11300 3445
rect 11370 3425 11390 3445
rect 11460 3425 11480 3445
rect 11550 3425 11570 3445
rect 11640 3425 11660 3445
rect 11730 3425 11750 3445
rect 11820 3425 11840 3445
rect 11910 3425 11930 3445
rect 12000 3425 12020 3445
rect 12090 3425 12110 3445
rect 12180 3425 12200 3445
rect 12270 3425 12290 3445
rect 12360 3425 12380 3445
rect 12450 3425 12470 3445
rect 12540 3425 12560 3445
rect 12630 3425 12650 3445
rect 12720 3425 12740 3445
rect 12810 3425 12830 3445
rect 12900 3425 12920 3445
rect 12990 3425 13010 3445
rect 13080 3425 13100 3445
rect 13170 3425 13190 3445
rect 13260 3425 13280 3445
rect 13350 3425 13370 3445
rect 13440 3425 13460 3445
rect 13530 3425 13550 3445
rect 13620 3425 13640 3445
rect 13710 3425 13730 3445
rect 13800 3425 13820 3445
rect 13890 3425 13910 3445
rect 13980 3425 14000 3445
rect 14070 3425 14090 3445
rect 14160 3425 14180 3445
rect 14250 3425 14270 3445
rect 14340 3425 14360 3445
rect 14430 3425 14450 3445
rect 14520 3425 14540 3445
rect 14610 3425 14630 3445
rect 14700 3425 14720 3445
rect 14790 3425 14810 3445
rect 14880 3425 14900 3445
rect 14970 3425 14990 3445
rect 15060 3425 15080 3445
rect 15150 3425 15170 3445
rect 15240 3425 15260 3445
rect 15330 3425 15350 3445
rect 15420 3425 15440 3445
rect 15510 3425 15530 3445
rect 15600 3425 15620 3445
rect 15690 3425 15710 3445
rect 15780 3425 15800 3445
rect 15870 3425 15890 3445
rect 15960 3425 15980 3445
rect 16050 3425 16070 3445
rect 16140 3425 16160 3445
rect 16230 3425 16250 3445
rect 16320 3425 16340 3445
rect 16410 3425 16430 3445
rect 16500 3425 16520 3445
rect 16590 3425 16610 3445
rect 16680 3425 16700 3445
rect 16770 3425 16790 3445
rect 16860 3425 16880 3445
rect 16950 3425 16970 3445
rect 17040 3425 17060 3445
rect 17130 3425 17150 3445
rect 17220 3425 17240 3445
rect 17310 3425 17330 3445
rect 17400 3425 17420 3445
rect 17490 3425 17510 3445
rect 17580 3425 17600 3445
rect 17670 3425 17690 3445
rect 17760 3425 17780 3445
rect 17850 3425 17870 3445
rect 17940 3425 17960 3445
rect 18030 3425 18050 3445
rect 18120 3425 18140 3445
rect 18210 3425 18230 3445
rect 18300 3425 18320 3445
rect 18390 3425 18410 3445
rect 18480 3425 18500 3445
rect 18570 3425 18590 3445
rect 18660 3425 18680 3445
rect 18750 3425 18770 3445
rect 18840 3425 18860 3445
rect 18930 3425 18950 3445
rect 19020 3425 19040 3445
rect 19110 3425 19130 3445
rect 19200 3425 19220 3445
rect 19290 3425 19310 3445
rect 19380 3425 19400 3445
rect 19470 3425 19490 3445
rect 19560 3425 19580 3445
rect 19650 3425 19670 3445
rect 19740 3425 19760 3445
rect 19830 3425 19850 3445
rect 19920 3425 19940 3445
rect 20010 3425 20030 3445
rect 20100 3425 20120 3445
rect 20190 3425 20210 3445
rect 20280 3425 20300 3445
rect 20370 3425 20390 3445
rect 20460 3425 20480 3445
rect 20550 3425 20570 3445
rect 20640 3425 20660 3445
<< nsubdiffcont >>
rect 9210 4345 9230 4365
rect 9300 4345 9320 4365
rect 9390 4345 9410 4365
rect 9480 4345 9500 4365
rect 9570 4345 9590 4365
rect 9660 4345 9680 4365
rect 9750 4345 9770 4365
rect 9840 4345 9860 4365
rect 9930 4345 9950 4365
rect 10020 4345 10040 4365
rect 10110 4345 10130 4365
rect 10200 4345 10220 4365
rect 10290 4345 10310 4365
rect 10380 4345 10400 4365
rect 10470 4345 10490 4365
rect 10560 4345 10580 4365
rect 10650 4345 10670 4365
rect 10740 4345 10760 4365
rect 10830 4345 10850 4365
rect 10920 4345 10940 4365
rect 11010 4345 11030 4365
rect 11100 4345 11120 4365
rect 11190 4345 11210 4365
rect 11280 4345 11300 4365
rect 11370 4345 11390 4365
rect 11460 4345 11480 4365
rect 11550 4345 11570 4365
rect 11640 4345 11660 4365
rect 11730 4345 11750 4365
rect 11820 4345 11840 4365
rect 11910 4345 11930 4365
rect 12000 4345 12020 4365
rect 12090 4345 12110 4365
rect 12180 4345 12200 4365
rect 12270 4345 12290 4365
rect 12360 4345 12380 4365
rect 12450 4345 12470 4365
rect 12540 4345 12560 4365
rect 12630 4345 12650 4365
rect 12720 4345 12740 4365
rect 12810 4345 12830 4365
rect 12900 4345 12920 4365
rect 12990 4345 13010 4365
rect 13080 4345 13100 4365
rect 13170 4345 13190 4365
rect 13260 4345 13280 4365
rect 13350 4345 13370 4365
rect 13440 4345 13460 4365
rect 13530 4345 13550 4365
rect 13620 4345 13640 4365
rect 13710 4345 13730 4365
rect 13800 4345 13820 4365
rect 13890 4345 13910 4365
rect 13980 4345 14000 4365
rect 14070 4345 14090 4365
rect 14160 4345 14180 4365
rect 14250 4345 14270 4365
rect 14340 4345 14360 4365
rect 14430 4345 14450 4365
rect 14520 4345 14540 4365
rect 14610 4345 14630 4365
rect 14700 4345 14720 4365
rect 14790 4345 14810 4365
rect 14880 4345 14900 4365
rect 14970 4345 14990 4365
rect 15060 4345 15080 4365
rect 15150 4345 15170 4365
rect 15240 4345 15260 4365
rect 15330 4345 15350 4365
rect 15420 4345 15440 4365
rect 15510 4345 15530 4365
rect 15600 4345 15620 4365
rect 15690 4345 15710 4365
rect 15780 4345 15800 4365
rect 15870 4345 15890 4365
rect 15960 4345 15980 4365
rect 16050 4345 16070 4365
rect 16140 4345 16160 4365
rect 16230 4345 16250 4365
rect 16320 4345 16340 4365
rect 16410 4345 16430 4365
rect 16500 4345 16520 4365
rect 16590 4345 16610 4365
rect 16680 4345 16700 4365
rect 16770 4345 16790 4365
rect 16860 4345 16880 4365
rect 16950 4345 16970 4365
rect 17040 4345 17060 4365
rect 17130 4345 17150 4365
rect 17220 4345 17240 4365
rect 17310 4345 17330 4365
rect 17400 4345 17420 4365
rect 17490 4345 17510 4365
rect 17580 4345 17600 4365
rect 17670 4345 17690 4365
rect 17760 4345 17780 4365
rect 17850 4345 17870 4365
rect 17940 4345 17960 4365
rect 18030 4345 18050 4365
rect 18120 4345 18140 4365
rect 18210 4345 18230 4365
rect 18300 4345 18320 4365
rect 18390 4345 18410 4365
rect 18480 4345 18500 4365
rect 18570 4345 18590 4365
rect 18660 4345 18680 4365
rect 18750 4345 18770 4365
rect 18840 4345 18860 4365
rect 18930 4345 18950 4365
rect 19020 4345 19040 4365
rect 19110 4345 19130 4365
rect 19200 4345 19220 4365
rect 19290 4345 19310 4365
rect 19380 4345 19400 4365
rect 19470 4345 19490 4365
rect 19560 4345 19580 4365
rect 19650 4345 19670 4365
rect 19740 4345 19760 4365
rect 19830 4345 19850 4365
rect 19920 4345 19940 4365
rect 20010 4345 20030 4365
rect 20100 4345 20120 4365
rect 20190 4345 20210 4365
rect 20280 4345 20300 4365
rect 20370 4345 20390 4365
rect 20460 4345 20480 4365
rect 20550 4345 20570 4365
rect 20640 4345 20660 4365
rect 9210 4125 9230 4145
rect 9300 4125 9320 4145
rect 9390 4125 9410 4145
rect 9480 4125 9500 4145
rect 9570 4125 9590 4145
rect 9660 4125 9680 4145
rect 9750 4125 9770 4145
rect 9840 4125 9860 4145
rect 9930 4125 9950 4145
rect 10020 4125 10040 4145
rect 10110 4125 10130 4145
rect 10200 4125 10220 4145
rect 10290 4125 10310 4145
rect 10380 4125 10400 4145
rect 10470 4125 10490 4145
rect 10560 4125 10580 4145
rect 10650 4125 10670 4145
rect 10740 4125 10760 4145
rect 10830 4125 10850 4145
rect 10920 4125 10940 4145
rect 11010 4125 11030 4145
rect 11100 4125 11120 4145
rect 11190 4125 11210 4145
rect 11280 4125 11300 4145
rect 11370 4125 11390 4145
rect 11460 4125 11480 4145
rect 11550 4125 11570 4145
rect 11640 4125 11660 4145
rect 11730 4125 11750 4145
rect 11820 4125 11840 4145
rect 11910 4125 11930 4145
rect 12000 4125 12020 4145
rect 12090 4125 12110 4145
rect 12180 4125 12200 4145
rect 12270 4125 12290 4145
rect 12360 4125 12380 4145
rect 12450 4125 12470 4145
rect 12540 4125 12560 4145
rect 12630 4125 12650 4145
rect 12720 4125 12740 4145
rect 12810 4125 12830 4145
rect 12900 4125 12920 4145
rect 12990 4125 13010 4145
rect 13080 4125 13100 4145
rect 13170 4125 13190 4145
rect 13260 4125 13280 4145
rect 13350 4125 13370 4145
rect 13440 4125 13460 4145
rect 13530 4125 13550 4145
rect 13620 4125 13640 4145
rect 13710 4125 13730 4145
rect 13800 4125 13820 4145
rect 13890 4125 13910 4145
rect 13980 4125 14000 4145
rect 14070 4125 14090 4145
rect 14160 4125 14180 4145
rect 14250 4125 14270 4145
rect 14340 4125 14360 4145
rect 14430 4125 14450 4145
rect 14520 4125 14540 4145
rect 14610 4125 14630 4145
rect 14700 4125 14720 4145
rect 14790 4125 14810 4145
rect 14880 4125 14900 4145
rect 14970 4125 14990 4145
rect 15060 4125 15080 4145
rect 15150 4125 15170 4145
rect 15240 4125 15260 4145
rect 15330 4125 15350 4145
rect 15420 4125 15440 4145
rect 15510 4125 15530 4145
rect 15600 4125 15620 4145
rect 15690 4125 15710 4145
rect 15780 4125 15800 4145
rect 15870 4125 15890 4145
rect 15960 4125 15980 4145
rect 16050 4125 16070 4145
rect 16140 4125 16160 4145
rect 16230 4125 16250 4145
rect 16320 4125 16340 4145
rect 16410 4125 16430 4145
rect 16500 4125 16520 4145
rect 16590 4125 16610 4145
rect 16680 4125 16700 4145
rect 16770 4125 16790 4145
rect 16860 4125 16880 4145
rect 16950 4125 16970 4145
rect 17040 4125 17060 4145
rect 17130 4125 17150 4145
rect 17220 4125 17240 4145
rect 17310 4125 17330 4145
rect 17400 4125 17420 4145
rect 17490 4125 17510 4145
rect 17580 4125 17600 4145
rect 17670 4125 17690 4145
rect 17760 4125 17780 4145
rect 17850 4125 17870 4145
rect 17940 4125 17960 4145
rect 18030 4125 18050 4145
rect 18120 4125 18140 4145
rect 18210 4125 18230 4145
rect 18300 4125 18320 4145
rect 18390 4125 18410 4145
rect 18480 4125 18500 4145
rect 18570 4125 18590 4145
rect 18660 4125 18680 4145
rect 18750 4125 18770 4145
rect 18840 4125 18860 4145
rect 18930 4125 18950 4145
rect 19020 4125 19040 4145
rect 19110 4125 19130 4145
rect 19200 4125 19220 4145
rect 19290 4125 19310 4145
rect 19380 4125 19400 4145
rect 19470 4125 19490 4145
rect 19560 4125 19580 4145
rect 19650 4125 19670 4145
rect 19740 4125 19760 4145
rect 19830 4125 19850 4145
rect 19920 4125 19940 4145
rect 20010 4125 20030 4145
rect 20100 4125 20120 4145
rect 20190 4125 20210 4145
rect 20280 4125 20300 4145
rect 20370 4125 20390 4145
rect 20460 4125 20480 4145
rect 20550 4125 20570 4145
rect 20640 4125 20660 4145
<< poly >>
rect 9195 4315 9245 4330
rect 9285 4315 9335 4330
rect 9375 4315 9425 4330
rect 9465 4315 9515 4330
rect 9555 4315 9605 4330
rect 9645 4315 9695 4330
rect 9735 4315 9785 4330
rect 9825 4315 9875 4330
rect 9915 4315 9965 4330
rect 10005 4315 10055 4330
rect 10095 4315 10145 4330
rect 10185 4315 10235 4330
rect 10275 4315 10325 4330
rect 10365 4315 10415 4330
rect 10455 4315 10505 4330
rect 10545 4315 10595 4330
rect 10635 4315 10685 4330
rect 10725 4315 10775 4330
rect 10815 4315 10865 4330
rect 10905 4315 10955 4330
rect 10995 4315 11045 4330
rect 11085 4315 11135 4330
rect 11175 4315 11225 4330
rect 11265 4315 11315 4330
rect 11355 4315 11405 4330
rect 11445 4315 11495 4330
rect 11535 4315 11585 4330
rect 11625 4315 11675 4330
rect 11715 4315 11765 4330
rect 11805 4315 11855 4330
rect 11895 4315 11945 4330
rect 11985 4315 12035 4330
rect 12075 4315 12125 4330
rect 12165 4315 12215 4330
rect 12255 4315 12305 4330
rect 12345 4315 12395 4330
rect 12435 4315 12485 4330
rect 12525 4315 12575 4330
rect 12615 4315 12665 4330
rect 12705 4315 12755 4330
rect 12795 4315 12845 4330
rect 12885 4315 12935 4330
rect 12975 4315 13025 4330
rect 13065 4315 13115 4330
rect 13155 4315 13205 4330
rect 13245 4315 13295 4330
rect 13335 4315 13385 4330
rect 13425 4315 13475 4330
rect 13515 4315 13565 4330
rect 13605 4315 13655 4330
rect 13695 4315 13745 4330
rect 13785 4315 13835 4330
rect 13875 4315 13925 4330
rect 13965 4315 14015 4330
rect 14055 4315 14105 4330
rect 14145 4315 14195 4330
rect 14235 4315 14285 4330
rect 14325 4315 14375 4330
rect 14415 4315 14465 4330
rect 14505 4315 14555 4330
rect 14595 4315 14645 4330
rect 14685 4315 14735 4330
rect 14775 4315 14825 4330
rect 14865 4315 14915 4330
rect 14955 4315 15005 4330
rect 15045 4315 15095 4330
rect 15135 4315 15185 4330
rect 15225 4315 15275 4330
rect 15315 4315 15365 4330
rect 15405 4315 15455 4330
rect 15495 4315 15545 4330
rect 15585 4315 15635 4330
rect 15675 4315 15725 4330
rect 15765 4315 15815 4330
rect 15855 4315 15905 4330
rect 15945 4315 15995 4330
rect 16035 4315 16085 4330
rect 16125 4315 16175 4330
rect 16215 4315 16265 4330
rect 16305 4315 16355 4330
rect 16395 4315 16445 4330
rect 16485 4315 16535 4330
rect 16575 4315 16625 4330
rect 16665 4315 16715 4330
rect 16755 4315 16805 4330
rect 16845 4315 16895 4330
rect 16935 4315 16985 4330
rect 17025 4315 17075 4330
rect 17115 4315 17165 4330
rect 17205 4315 17255 4330
rect 17295 4315 17345 4330
rect 17385 4315 17435 4330
rect 17475 4315 17525 4330
rect 17565 4315 17615 4330
rect 17655 4315 17705 4330
rect 17745 4315 17795 4330
rect 17835 4315 17885 4330
rect 17925 4315 17975 4330
rect 18015 4315 18065 4330
rect 18105 4315 18155 4330
rect 18195 4315 18245 4330
rect 18285 4315 18335 4330
rect 18375 4315 18425 4330
rect 18465 4315 18515 4330
rect 18555 4315 18605 4330
rect 18645 4315 18695 4330
rect 18735 4315 18785 4330
rect 18825 4315 18875 4330
rect 18915 4315 18965 4330
rect 19005 4315 19055 4330
rect 19095 4315 19145 4330
rect 19185 4315 19235 4330
rect 19275 4315 19325 4330
rect 19365 4315 19415 4330
rect 19455 4315 19505 4330
rect 19545 4315 19595 4330
rect 19635 4315 19685 4330
rect 19725 4315 19775 4330
rect 19815 4315 19865 4330
rect 19905 4315 19955 4330
rect 19995 4315 20045 4330
rect 20085 4315 20135 4330
rect 20175 4315 20225 4330
rect 20265 4315 20315 4330
rect 20355 4315 20405 4330
rect 20445 4315 20495 4330
rect 20535 4315 20585 4330
rect 20625 4315 20675 4330
rect 9195 4195 9245 4215
rect 9285 4195 9335 4215
rect 9195 4190 9335 4195
rect 9195 4170 9210 4190
rect 9230 4170 9300 4190
rect 9320 4170 9335 4190
rect 9195 4165 9335 4170
rect 9375 4195 9425 4215
rect 9465 4195 9515 4215
rect 9375 4190 9515 4195
rect 9375 4170 9390 4190
rect 9410 4170 9480 4190
rect 9500 4170 9515 4190
rect 9375 4165 9515 4170
rect 9555 4195 9605 4215
rect 9645 4195 9695 4215
rect 9555 4190 9695 4195
rect 9555 4170 9570 4190
rect 9590 4170 9660 4190
rect 9680 4170 9695 4190
rect 9555 4165 9695 4170
rect 9735 4195 9785 4215
rect 9825 4195 9875 4215
rect 9735 4190 9875 4195
rect 9735 4170 9750 4190
rect 9770 4170 9840 4190
rect 9860 4170 9875 4190
rect 9735 4165 9875 4170
rect 9915 4195 9965 4215
rect 10005 4195 10055 4215
rect 9915 4190 10055 4195
rect 9915 4170 9930 4190
rect 9950 4170 10020 4190
rect 10040 4170 10055 4190
rect 9915 4165 10055 4170
rect 10095 4195 10145 4215
rect 10185 4195 10235 4215
rect 10095 4190 10235 4195
rect 10095 4170 10110 4190
rect 10130 4170 10200 4190
rect 10220 4170 10235 4190
rect 10095 4165 10235 4170
rect 10275 4195 10325 4215
rect 10365 4195 10415 4215
rect 10275 4190 10415 4195
rect 10275 4170 10290 4190
rect 10310 4170 10380 4190
rect 10400 4170 10415 4190
rect 10275 4165 10415 4170
rect 10455 4195 10505 4215
rect 10545 4195 10595 4215
rect 10455 4190 10595 4195
rect 10455 4170 10470 4190
rect 10490 4170 10560 4190
rect 10580 4170 10595 4190
rect 10455 4165 10595 4170
rect 10635 4195 10685 4215
rect 10725 4195 10775 4215
rect 10635 4190 10775 4195
rect 10635 4170 10650 4190
rect 10670 4170 10740 4190
rect 10760 4170 10775 4190
rect 10635 4165 10775 4170
rect 10815 4195 10865 4215
rect 10905 4195 10955 4215
rect 10815 4190 10955 4195
rect 10815 4170 10830 4190
rect 10850 4170 10920 4190
rect 10940 4170 10955 4190
rect 10815 4165 10955 4170
rect 10995 4195 11045 4215
rect 11085 4195 11135 4215
rect 10995 4190 11135 4195
rect 10995 4170 11010 4190
rect 11030 4170 11100 4190
rect 11120 4170 11135 4190
rect 10995 4165 11135 4170
rect 11175 4195 11225 4215
rect 11265 4195 11315 4215
rect 11175 4190 11315 4195
rect 11175 4170 11190 4190
rect 11210 4170 11280 4190
rect 11300 4170 11315 4190
rect 11175 4165 11315 4170
rect 11355 4195 11405 4215
rect 11445 4195 11495 4215
rect 11355 4190 11495 4195
rect 11355 4170 11370 4190
rect 11390 4170 11460 4190
rect 11480 4170 11495 4190
rect 11355 4165 11495 4170
rect 11535 4195 11585 4215
rect 11625 4195 11675 4215
rect 11535 4190 11675 4195
rect 11535 4170 11550 4190
rect 11570 4170 11640 4190
rect 11660 4170 11675 4190
rect 11535 4165 11675 4170
rect 11715 4195 11765 4215
rect 11805 4195 11855 4215
rect 11715 4190 11855 4195
rect 11715 4170 11730 4190
rect 11750 4170 11820 4190
rect 11840 4170 11855 4190
rect 11715 4165 11855 4170
rect 11895 4195 11945 4215
rect 11985 4195 12035 4215
rect 11895 4190 12035 4195
rect 11895 4170 11910 4190
rect 11930 4170 12000 4190
rect 12020 4170 12035 4190
rect 11895 4165 12035 4170
rect 12075 4195 12125 4215
rect 12165 4195 12215 4215
rect 12075 4190 12215 4195
rect 12075 4170 12090 4190
rect 12110 4170 12180 4190
rect 12200 4170 12215 4190
rect 12075 4165 12215 4170
rect 12255 4195 12305 4215
rect 12345 4195 12395 4215
rect 12255 4190 12395 4195
rect 12255 4170 12270 4190
rect 12290 4170 12360 4190
rect 12380 4170 12395 4190
rect 12255 4165 12395 4170
rect 12435 4195 12485 4215
rect 12525 4195 12575 4215
rect 12435 4190 12575 4195
rect 12435 4170 12450 4190
rect 12470 4170 12540 4190
rect 12560 4170 12575 4190
rect 12435 4165 12575 4170
rect 12615 4195 12665 4215
rect 12705 4195 12755 4215
rect 12615 4190 12755 4195
rect 12615 4170 12630 4190
rect 12650 4170 12720 4190
rect 12740 4170 12755 4190
rect 12615 4165 12755 4170
rect 12795 4195 12845 4215
rect 12885 4195 12935 4215
rect 12795 4190 12935 4195
rect 12795 4170 12810 4190
rect 12830 4170 12900 4190
rect 12920 4170 12935 4190
rect 12795 4165 12935 4170
rect 12975 4195 13025 4215
rect 13065 4195 13115 4215
rect 12975 4190 13115 4195
rect 12975 4170 12990 4190
rect 13010 4170 13080 4190
rect 13100 4170 13115 4190
rect 12975 4165 13115 4170
rect 13155 4195 13205 4215
rect 13245 4195 13295 4215
rect 13155 4190 13295 4195
rect 13155 4170 13170 4190
rect 13190 4170 13260 4190
rect 13280 4170 13295 4190
rect 13155 4165 13295 4170
rect 13335 4195 13385 4215
rect 13425 4195 13475 4215
rect 13335 4190 13475 4195
rect 13335 4170 13350 4190
rect 13370 4170 13440 4190
rect 13460 4170 13475 4190
rect 13335 4165 13475 4170
rect 13515 4195 13565 4215
rect 13605 4195 13655 4215
rect 13515 4190 13655 4195
rect 13515 4170 13530 4190
rect 13550 4170 13620 4190
rect 13640 4170 13655 4190
rect 13515 4165 13655 4170
rect 13695 4195 13745 4215
rect 13785 4195 13835 4215
rect 13695 4190 13835 4195
rect 13695 4170 13710 4190
rect 13730 4170 13800 4190
rect 13820 4170 13835 4190
rect 13695 4165 13835 4170
rect 13875 4195 13925 4215
rect 13965 4195 14015 4215
rect 13875 4190 14015 4195
rect 13875 4170 13890 4190
rect 13910 4170 13980 4190
rect 14000 4170 14015 4190
rect 13875 4165 14015 4170
rect 14055 4195 14105 4215
rect 14145 4195 14195 4215
rect 14055 4190 14195 4195
rect 14055 4170 14070 4190
rect 14090 4170 14160 4190
rect 14180 4170 14195 4190
rect 14055 4165 14195 4170
rect 14235 4195 14285 4215
rect 14325 4195 14375 4215
rect 14235 4190 14375 4195
rect 14235 4170 14250 4190
rect 14270 4170 14340 4190
rect 14360 4170 14375 4190
rect 14235 4165 14375 4170
rect 14415 4195 14465 4215
rect 14505 4195 14555 4215
rect 14415 4190 14555 4195
rect 14415 4170 14430 4190
rect 14450 4170 14520 4190
rect 14540 4170 14555 4190
rect 14415 4165 14555 4170
rect 14595 4195 14645 4215
rect 14685 4195 14735 4215
rect 14595 4190 14735 4195
rect 14595 4170 14610 4190
rect 14630 4170 14700 4190
rect 14720 4170 14735 4190
rect 14595 4165 14735 4170
rect 14775 4195 14825 4215
rect 14865 4195 14915 4215
rect 14775 4190 14915 4195
rect 14775 4170 14790 4190
rect 14810 4170 14880 4190
rect 14900 4170 14915 4190
rect 14775 4165 14915 4170
rect 14955 4195 15005 4215
rect 15045 4195 15095 4215
rect 14955 4190 15095 4195
rect 14955 4170 14970 4190
rect 14990 4170 15060 4190
rect 15080 4170 15095 4190
rect 14955 4165 15095 4170
rect 15135 4195 15185 4215
rect 15225 4195 15275 4215
rect 15135 4190 15275 4195
rect 15135 4170 15150 4190
rect 15170 4170 15240 4190
rect 15260 4170 15275 4190
rect 15135 4165 15275 4170
rect 15315 4195 15365 4215
rect 15405 4195 15455 4215
rect 15315 4190 15455 4195
rect 15315 4170 15330 4190
rect 15350 4170 15420 4190
rect 15440 4170 15455 4190
rect 15315 4165 15455 4170
rect 15495 4195 15545 4215
rect 15585 4195 15635 4215
rect 15495 4190 15635 4195
rect 15495 4170 15510 4190
rect 15530 4170 15600 4190
rect 15620 4170 15635 4190
rect 15495 4165 15635 4170
rect 15675 4195 15725 4215
rect 15765 4195 15815 4215
rect 15675 4190 15815 4195
rect 15675 4170 15690 4190
rect 15710 4170 15780 4190
rect 15800 4170 15815 4190
rect 15675 4165 15815 4170
rect 15855 4195 15905 4215
rect 15945 4195 15995 4215
rect 15855 4190 15995 4195
rect 15855 4170 15870 4190
rect 15890 4170 15960 4190
rect 15980 4170 15995 4190
rect 15855 4165 15995 4170
rect 16035 4195 16085 4215
rect 16125 4195 16175 4215
rect 16035 4190 16175 4195
rect 16035 4170 16050 4190
rect 16070 4170 16140 4190
rect 16160 4170 16175 4190
rect 16035 4165 16175 4170
rect 16215 4195 16265 4215
rect 16305 4195 16355 4215
rect 16215 4190 16355 4195
rect 16215 4170 16230 4190
rect 16250 4170 16320 4190
rect 16340 4170 16355 4190
rect 16215 4165 16355 4170
rect 16395 4195 16445 4215
rect 16485 4195 16535 4215
rect 16395 4190 16535 4195
rect 16395 4170 16410 4190
rect 16430 4170 16500 4190
rect 16520 4170 16535 4190
rect 16395 4165 16535 4170
rect 16575 4195 16625 4215
rect 16665 4195 16715 4215
rect 16575 4190 16715 4195
rect 16575 4170 16590 4190
rect 16610 4170 16680 4190
rect 16700 4170 16715 4190
rect 16575 4165 16715 4170
rect 16755 4195 16805 4215
rect 16845 4195 16895 4215
rect 16755 4190 16895 4195
rect 16755 4170 16770 4190
rect 16790 4170 16860 4190
rect 16880 4170 16895 4190
rect 16755 4165 16895 4170
rect 16935 4195 16985 4215
rect 17025 4195 17075 4215
rect 16935 4190 17075 4195
rect 16935 4170 16950 4190
rect 16970 4170 17040 4190
rect 17060 4170 17075 4190
rect 16935 4165 17075 4170
rect 17115 4195 17165 4215
rect 17205 4195 17255 4215
rect 17115 4190 17255 4195
rect 17115 4170 17130 4190
rect 17150 4170 17220 4190
rect 17240 4170 17255 4190
rect 17115 4165 17255 4170
rect 17295 4195 17345 4215
rect 17385 4195 17435 4215
rect 17295 4190 17435 4195
rect 17295 4170 17310 4190
rect 17330 4170 17400 4190
rect 17420 4170 17435 4190
rect 17295 4165 17435 4170
rect 17475 4195 17525 4215
rect 17565 4195 17615 4215
rect 17475 4190 17615 4195
rect 17475 4170 17490 4190
rect 17510 4170 17580 4190
rect 17600 4170 17615 4190
rect 17475 4165 17615 4170
rect 17655 4195 17705 4215
rect 17745 4195 17795 4215
rect 17655 4190 17795 4195
rect 17655 4170 17670 4190
rect 17690 4170 17760 4190
rect 17780 4170 17795 4190
rect 17655 4165 17795 4170
rect 17835 4195 17885 4215
rect 17925 4195 17975 4215
rect 17835 4190 17975 4195
rect 17835 4170 17850 4190
rect 17870 4170 17940 4190
rect 17960 4170 17975 4190
rect 17835 4165 17975 4170
rect 18015 4195 18065 4215
rect 18105 4195 18155 4215
rect 18015 4190 18155 4195
rect 18015 4170 18030 4190
rect 18050 4170 18120 4190
rect 18140 4170 18155 4190
rect 18015 4165 18155 4170
rect 18195 4195 18245 4215
rect 18285 4195 18335 4215
rect 18195 4190 18335 4195
rect 18195 4170 18210 4190
rect 18230 4170 18300 4190
rect 18320 4170 18335 4190
rect 18195 4165 18335 4170
rect 18375 4195 18425 4215
rect 18465 4195 18515 4215
rect 18375 4190 18515 4195
rect 18375 4170 18390 4190
rect 18410 4170 18480 4190
rect 18500 4170 18515 4190
rect 18375 4165 18515 4170
rect 18555 4195 18605 4215
rect 18645 4195 18695 4215
rect 18555 4190 18695 4195
rect 18555 4170 18570 4190
rect 18590 4170 18660 4190
rect 18680 4170 18695 4190
rect 18555 4165 18695 4170
rect 18735 4195 18785 4215
rect 18825 4195 18875 4215
rect 18735 4190 18875 4195
rect 18735 4170 18750 4190
rect 18770 4170 18840 4190
rect 18860 4170 18875 4190
rect 18735 4165 18875 4170
rect 18915 4195 18965 4215
rect 19005 4195 19055 4215
rect 18915 4190 19055 4195
rect 18915 4170 18930 4190
rect 18950 4170 19020 4190
rect 19040 4170 19055 4190
rect 18915 4165 19055 4170
rect 19095 4195 19145 4215
rect 19185 4195 19235 4215
rect 19095 4190 19235 4195
rect 19095 4170 19110 4190
rect 19130 4170 19200 4190
rect 19220 4170 19235 4190
rect 19095 4165 19235 4170
rect 19275 4195 19325 4215
rect 19365 4195 19415 4215
rect 19275 4190 19415 4195
rect 19275 4170 19290 4190
rect 19310 4170 19380 4190
rect 19400 4170 19415 4190
rect 19275 4165 19415 4170
rect 19455 4195 19505 4215
rect 19545 4195 19595 4215
rect 19455 4190 19595 4195
rect 19455 4170 19470 4190
rect 19490 4170 19560 4190
rect 19580 4170 19595 4190
rect 19455 4165 19595 4170
rect 19635 4195 19685 4215
rect 19725 4195 19775 4215
rect 19635 4190 19775 4195
rect 19635 4170 19650 4190
rect 19670 4170 19740 4190
rect 19760 4170 19775 4190
rect 19635 4165 19775 4170
rect 19815 4195 19865 4215
rect 19905 4195 19955 4215
rect 19815 4190 19955 4195
rect 19815 4170 19830 4190
rect 19850 4170 19920 4190
rect 19940 4170 19955 4190
rect 19815 4165 19955 4170
rect 19995 4195 20045 4215
rect 20085 4195 20135 4215
rect 19995 4190 20135 4195
rect 19995 4170 20010 4190
rect 20030 4170 20100 4190
rect 20120 4170 20135 4190
rect 19995 4165 20135 4170
rect 20175 4195 20225 4215
rect 20265 4195 20315 4215
rect 20175 4190 20315 4195
rect 20175 4170 20190 4190
rect 20210 4170 20280 4190
rect 20300 4170 20315 4190
rect 20175 4165 20315 4170
rect 20355 4195 20405 4215
rect 20445 4195 20495 4215
rect 20355 4190 20495 4195
rect 20355 4170 20370 4190
rect 20390 4170 20460 4190
rect 20480 4170 20495 4190
rect 20355 4165 20495 4170
rect 20535 4195 20585 4215
rect 20625 4195 20675 4215
rect 20535 4190 20675 4195
rect 20535 4170 20550 4190
rect 20570 4170 20640 4190
rect 20660 4170 20675 4190
rect 20535 4165 20675 4170
rect 9195 3620 9335 3625
rect 9195 3600 9210 3620
rect 9230 3600 9300 3620
rect 9320 3600 9335 3620
rect 9195 3595 9335 3600
rect 9195 3575 9245 3595
rect 9285 3575 9335 3595
rect 9375 3620 9515 3625
rect 9375 3600 9390 3620
rect 9410 3600 9480 3620
rect 9500 3600 9515 3620
rect 9375 3595 9515 3600
rect 9375 3575 9425 3595
rect 9465 3575 9515 3595
rect 9555 3620 9695 3625
rect 9555 3600 9570 3620
rect 9590 3600 9660 3620
rect 9680 3600 9695 3620
rect 9555 3595 9695 3600
rect 9555 3575 9605 3595
rect 9645 3575 9695 3595
rect 9735 3620 9875 3625
rect 9735 3600 9750 3620
rect 9770 3600 9840 3620
rect 9860 3600 9875 3620
rect 9735 3595 9875 3600
rect 9735 3575 9785 3595
rect 9825 3575 9875 3595
rect 9915 3620 10055 3625
rect 9915 3600 9930 3620
rect 9950 3600 10020 3620
rect 10040 3600 10055 3620
rect 9915 3595 10055 3600
rect 9915 3575 9965 3595
rect 10005 3575 10055 3595
rect 10095 3620 10235 3625
rect 10095 3600 10110 3620
rect 10130 3600 10200 3620
rect 10220 3600 10235 3620
rect 10095 3595 10235 3600
rect 10095 3575 10145 3595
rect 10185 3575 10235 3595
rect 10275 3620 10415 3625
rect 10275 3600 10290 3620
rect 10310 3600 10380 3620
rect 10400 3600 10415 3620
rect 10275 3595 10415 3600
rect 10275 3575 10325 3595
rect 10365 3575 10415 3595
rect 10455 3620 10595 3625
rect 10455 3600 10470 3620
rect 10490 3600 10560 3620
rect 10580 3600 10595 3620
rect 10455 3595 10595 3600
rect 10455 3575 10505 3595
rect 10545 3575 10595 3595
rect 10635 3620 10775 3625
rect 10635 3600 10650 3620
rect 10670 3600 10740 3620
rect 10760 3600 10775 3620
rect 10635 3595 10775 3600
rect 10635 3575 10685 3595
rect 10725 3575 10775 3595
rect 10815 3620 10955 3625
rect 10815 3600 10830 3620
rect 10850 3600 10920 3620
rect 10940 3600 10955 3620
rect 10815 3595 10955 3600
rect 10815 3575 10865 3595
rect 10905 3575 10955 3595
rect 10995 3620 11135 3625
rect 10995 3600 11010 3620
rect 11030 3600 11100 3620
rect 11120 3600 11135 3620
rect 10995 3595 11135 3600
rect 10995 3575 11045 3595
rect 11085 3575 11135 3595
rect 11175 3620 11315 3625
rect 11175 3600 11190 3620
rect 11210 3600 11280 3620
rect 11300 3600 11315 3620
rect 11175 3595 11315 3600
rect 11175 3575 11225 3595
rect 11265 3575 11315 3595
rect 11355 3620 11495 3625
rect 11355 3600 11370 3620
rect 11390 3600 11460 3620
rect 11480 3600 11495 3620
rect 11355 3595 11495 3600
rect 11355 3575 11405 3595
rect 11445 3575 11495 3595
rect 11535 3620 11675 3625
rect 11535 3600 11550 3620
rect 11570 3600 11640 3620
rect 11660 3600 11675 3620
rect 11535 3595 11675 3600
rect 11535 3575 11585 3595
rect 11625 3575 11675 3595
rect 11715 3620 11855 3625
rect 11715 3600 11730 3620
rect 11750 3600 11820 3620
rect 11840 3600 11855 3620
rect 11715 3595 11855 3600
rect 11715 3575 11765 3595
rect 11805 3575 11855 3595
rect 11895 3620 12035 3625
rect 11895 3600 11910 3620
rect 11930 3600 12000 3620
rect 12020 3600 12035 3620
rect 11895 3595 12035 3600
rect 11895 3575 11945 3595
rect 11985 3575 12035 3595
rect 12075 3620 12215 3625
rect 12075 3600 12090 3620
rect 12110 3600 12180 3620
rect 12200 3600 12215 3620
rect 12075 3595 12215 3600
rect 12075 3575 12125 3595
rect 12165 3575 12215 3595
rect 12255 3620 12395 3625
rect 12255 3600 12270 3620
rect 12290 3600 12360 3620
rect 12380 3600 12395 3620
rect 12255 3595 12395 3600
rect 12255 3575 12305 3595
rect 12345 3575 12395 3595
rect 12435 3620 12575 3625
rect 12435 3600 12450 3620
rect 12470 3600 12540 3620
rect 12560 3600 12575 3620
rect 12435 3595 12575 3600
rect 12435 3575 12485 3595
rect 12525 3575 12575 3595
rect 12615 3620 12755 3625
rect 12615 3600 12630 3620
rect 12650 3600 12720 3620
rect 12740 3600 12755 3620
rect 12615 3595 12755 3600
rect 12615 3575 12665 3595
rect 12705 3575 12755 3595
rect 12795 3620 12935 3625
rect 12795 3600 12810 3620
rect 12830 3600 12900 3620
rect 12920 3600 12935 3620
rect 12795 3595 12935 3600
rect 12795 3575 12845 3595
rect 12885 3575 12935 3595
rect 12975 3620 13115 3625
rect 12975 3600 12990 3620
rect 13010 3600 13080 3620
rect 13100 3600 13115 3620
rect 12975 3595 13115 3600
rect 12975 3575 13025 3595
rect 13065 3575 13115 3595
rect 13155 3620 13295 3625
rect 13155 3600 13170 3620
rect 13190 3600 13260 3620
rect 13280 3600 13295 3620
rect 13155 3595 13295 3600
rect 13155 3575 13205 3595
rect 13245 3575 13295 3595
rect 13335 3620 13475 3625
rect 13335 3600 13350 3620
rect 13370 3600 13440 3620
rect 13460 3600 13475 3620
rect 13335 3595 13475 3600
rect 13335 3575 13385 3595
rect 13425 3575 13475 3595
rect 13515 3620 13655 3625
rect 13515 3600 13530 3620
rect 13550 3600 13620 3620
rect 13640 3600 13655 3620
rect 13515 3595 13655 3600
rect 13515 3575 13565 3595
rect 13605 3575 13655 3595
rect 13695 3620 13835 3625
rect 13695 3600 13710 3620
rect 13730 3600 13800 3620
rect 13820 3600 13835 3620
rect 13695 3595 13835 3600
rect 13695 3575 13745 3595
rect 13785 3575 13835 3595
rect 13875 3620 14015 3625
rect 13875 3600 13890 3620
rect 13910 3600 13980 3620
rect 14000 3600 14015 3620
rect 13875 3595 14015 3600
rect 13875 3575 13925 3595
rect 13965 3575 14015 3595
rect 14055 3620 14195 3625
rect 14055 3600 14070 3620
rect 14090 3600 14160 3620
rect 14180 3600 14195 3620
rect 14055 3595 14195 3600
rect 14055 3575 14105 3595
rect 14145 3575 14195 3595
rect 14235 3620 14375 3625
rect 14235 3600 14250 3620
rect 14270 3600 14340 3620
rect 14360 3600 14375 3620
rect 14235 3595 14375 3600
rect 14235 3575 14285 3595
rect 14325 3575 14375 3595
rect 14415 3620 14555 3625
rect 14415 3600 14430 3620
rect 14450 3600 14520 3620
rect 14540 3600 14555 3620
rect 14415 3595 14555 3600
rect 14415 3575 14465 3595
rect 14505 3575 14555 3595
rect 14595 3620 14735 3625
rect 14595 3600 14610 3620
rect 14630 3600 14700 3620
rect 14720 3600 14735 3620
rect 14595 3595 14735 3600
rect 14595 3575 14645 3595
rect 14685 3575 14735 3595
rect 14775 3620 14915 3625
rect 14775 3600 14790 3620
rect 14810 3600 14880 3620
rect 14900 3600 14915 3620
rect 14775 3595 14915 3600
rect 14775 3575 14825 3595
rect 14865 3575 14915 3595
rect 14955 3620 15095 3625
rect 14955 3600 14970 3620
rect 14990 3600 15060 3620
rect 15080 3600 15095 3620
rect 14955 3595 15095 3600
rect 14955 3575 15005 3595
rect 15045 3575 15095 3595
rect 15135 3620 15275 3625
rect 15135 3600 15150 3620
rect 15170 3600 15240 3620
rect 15260 3600 15275 3620
rect 15135 3595 15275 3600
rect 15135 3575 15185 3595
rect 15225 3575 15275 3595
rect 15315 3620 15455 3625
rect 15315 3600 15330 3620
rect 15350 3600 15420 3620
rect 15440 3600 15455 3620
rect 15315 3595 15455 3600
rect 15315 3575 15365 3595
rect 15405 3575 15455 3595
rect 15495 3620 15635 3625
rect 15495 3600 15510 3620
rect 15530 3600 15600 3620
rect 15620 3600 15635 3620
rect 15495 3595 15635 3600
rect 15495 3575 15545 3595
rect 15585 3575 15635 3595
rect 15675 3620 15815 3625
rect 15675 3600 15690 3620
rect 15710 3600 15780 3620
rect 15800 3600 15815 3620
rect 15675 3595 15815 3600
rect 15675 3575 15725 3595
rect 15765 3575 15815 3595
rect 15855 3620 15995 3625
rect 15855 3600 15870 3620
rect 15890 3600 15960 3620
rect 15980 3600 15995 3620
rect 15855 3595 15995 3600
rect 15855 3575 15905 3595
rect 15945 3575 15995 3595
rect 16035 3620 16175 3625
rect 16035 3600 16050 3620
rect 16070 3600 16140 3620
rect 16160 3600 16175 3620
rect 16035 3595 16175 3600
rect 16035 3575 16085 3595
rect 16125 3575 16175 3595
rect 16215 3620 16355 3625
rect 16215 3600 16230 3620
rect 16250 3600 16320 3620
rect 16340 3600 16355 3620
rect 16215 3595 16355 3600
rect 16215 3575 16265 3595
rect 16305 3575 16355 3595
rect 16395 3620 16535 3625
rect 16395 3600 16410 3620
rect 16430 3600 16500 3620
rect 16520 3600 16535 3620
rect 16395 3595 16535 3600
rect 16395 3575 16445 3595
rect 16485 3575 16535 3595
rect 16575 3620 16715 3625
rect 16575 3600 16590 3620
rect 16610 3600 16680 3620
rect 16700 3600 16715 3620
rect 16575 3595 16715 3600
rect 16575 3575 16625 3595
rect 16665 3575 16715 3595
rect 16755 3620 16895 3625
rect 16755 3600 16770 3620
rect 16790 3600 16860 3620
rect 16880 3600 16895 3620
rect 16755 3595 16895 3600
rect 16755 3575 16805 3595
rect 16845 3575 16895 3595
rect 16935 3620 17075 3625
rect 16935 3600 16950 3620
rect 16970 3600 17040 3620
rect 17060 3600 17075 3620
rect 16935 3595 17075 3600
rect 16935 3575 16985 3595
rect 17025 3575 17075 3595
rect 17115 3620 17255 3625
rect 17115 3600 17130 3620
rect 17150 3600 17220 3620
rect 17240 3600 17255 3620
rect 17115 3595 17255 3600
rect 17115 3575 17165 3595
rect 17205 3575 17255 3595
rect 17295 3620 17435 3625
rect 17295 3600 17310 3620
rect 17330 3600 17400 3620
rect 17420 3600 17435 3620
rect 17295 3595 17435 3600
rect 17295 3575 17345 3595
rect 17385 3575 17435 3595
rect 17475 3620 17615 3625
rect 17475 3600 17490 3620
rect 17510 3600 17580 3620
rect 17600 3600 17615 3620
rect 17475 3595 17615 3600
rect 17475 3575 17525 3595
rect 17565 3575 17615 3595
rect 17655 3620 17795 3625
rect 17655 3600 17670 3620
rect 17690 3600 17760 3620
rect 17780 3600 17795 3620
rect 17655 3595 17795 3600
rect 17655 3575 17705 3595
rect 17745 3575 17795 3595
rect 17835 3620 17975 3625
rect 17835 3600 17850 3620
rect 17870 3600 17940 3620
rect 17960 3600 17975 3620
rect 17835 3595 17975 3600
rect 17835 3575 17885 3595
rect 17925 3575 17975 3595
rect 18015 3620 18155 3625
rect 18015 3600 18030 3620
rect 18050 3600 18120 3620
rect 18140 3600 18155 3620
rect 18015 3595 18155 3600
rect 18015 3575 18065 3595
rect 18105 3575 18155 3595
rect 18195 3620 18335 3625
rect 18195 3600 18210 3620
rect 18230 3600 18300 3620
rect 18320 3600 18335 3620
rect 18195 3595 18335 3600
rect 18195 3575 18245 3595
rect 18285 3575 18335 3595
rect 18375 3620 18515 3625
rect 18375 3600 18390 3620
rect 18410 3600 18480 3620
rect 18500 3600 18515 3620
rect 18375 3595 18515 3600
rect 18375 3575 18425 3595
rect 18465 3575 18515 3595
rect 18555 3620 18695 3625
rect 18555 3600 18570 3620
rect 18590 3600 18660 3620
rect 18680 3600 18695 3620
rect 18555 3595 18695 3600
rect 18555 3575 18605 3595
rect 18645 3575 18695 3595
rect 18735 3620 18875 3625
rect 18735 3600 18750 3620
rect 18770 3600 18840 3620
rect 18860 3600 18875 3620
rect 18735 3595 18875 3600
rect 18735 3575 18785 3595
rect 18825 3575 18875 3595
rect 18915 3620 19055 3625
rect 18915 3600 18930 3620
rect 18950 3600 19020 3620
rect 19040 3600 19055 3620
rect 18915 3595 19055 3600
rect 18915 3575 18965 3595
rect 19005 3575 19055 3595
rect 19095 3620 19235 3625
rect 19095 3600 19110 3620
rect 19130 3600 19200 3620
rect 19220 3600 19235 3620
rect 19095 3595 19235 3600
rect 19095 3575 19145 3595
rect 19185 3575 19235 3595
rect 19275 3620 19415 3625
rect 19275 3600 19290 3620
rect 19310 3600 19380 3620
rect 19400 3600 19415 3620
rect 19275 3595 19415 3600
rect 19275 3575 19325 3595
rect 19365 3575 19415 3595
rect 19455 3620 19595 3625
rect 19455 3600 19470 3620
rect 19490 3600 19560 3620
rect 19580 3600 19595 3620
rect 19455 3595 19595 3600
rect 19455 3575 19505 3595
rect 19545 3575 19595 3595
rect 19635 3620 19775 3625
rect 19635 3600 19650 3620
rect 19670 3600 19740 3620
rect 19760 3600 19775 3620
rect 19635 3595 19775 3600
rect 19635 3575 19685 3595
rect 19725 3575 19775 3595
rect 19815 3620 19955 3625
rect 19815 3600 19830 3620
rect 19850 3600 19920 3620
rect 19940 3600 19955 3620
rect 19815 3595 19955 3600
rect 19815 3575 19865 3595
rect 19905 3575 19955 3595
rect 19995 3620 20135 3625
rect 19995 3600 20010 3620
rect 20030 3600 20100 3620
rect 20120 3600 20135 3620
rect 19995 3595 20135 3600
rect 19995 3575 20045 3595
rect 20085 3575 20135 3595
rect 20175 3620 20315 3625
rect 20175 3600 20190 3620
rect 20210 3600 20280 3620
rect 20300 3600 20315 3620
rect 20175 3595 20315 3600
rect 20175 3575 20225 3595
rect 20265 3575 20315 3595
rect 20355 3620 20495 3625
rect 20355 3600 20370 3620
rect 20390 3600 20460 3620
rect 20480 3600 20495 3620
rect 20355 3595 20495 3600
rect 20355 3575 20405 3595
rect 20445 3575 20495 3595
rect 20535 3620 20675 3625
rect 20535 3600 20550 3620
rect 20570 3600 20640 3620
rect 20660 3600 20675 3620
rect 20535 3595 20675 3600
rect 20535 3575 20585 3595
rect 20625 3575 20675 3595
rect 9195 3460 9245 3475
rect 9285 3460 9335 3475
rect 9375 3460 9425 3475
rect 9465 3460 9515 3475
rect 9555 3460 9605 3475
rect 9645 3460 9695 3475
rect 9735 3460 9785 3475
rect 9825 3460 9875 3475
rect 9915 3460 9965 3475
rect 10005 3460 10055 3475
rect 10095 3460 10145 3475
rect 10185 3460 10235 3475
rect 10275 3460 10325 3475
rect 10365 3460 10415 3475
rect 10455 3460 10505 3475
rect 10545 3460 10595 3475
rect 10635 3460 10685 3475
rect 10725 3460 10775 3475
rect 10815 3460 10865 3475
rect 10905 3460 10955 3475
rect 10995 3460 11045 3475
rect 11085 3460 11135 3475
rect 11175 3460 11225 3475
rect 11265 3460 11315 3475
rect 11355 3460 11405 3475
rect 11445 3460 11495 3475
rect 11535 3460 11585 3475
rect 11625 3460 11675 3475
rect 11715 3460 11765 3475
rect 11805 3460 11855 3475
rect 11895 3460 11945 3475
rect 11985 3460 12035 3475
rect 12075 3460 12125 3475
rect 12165 3460 12215 3475
rect 12255 3460 12305 3475
rect 12345 3460 12395 3475
rect 12435 3460 12485 3475
rect 12525 3460 12575 3475
rect 12615 3460 12665 3475
rect 12705 3460 12755 3475
rect 12795 3460 12845 3475
rect 12885 3460 12935 3475
rect 12975 3460 13025 3475
rect 13065 3460 13115 3475
rect 13155 3460 13205 3475
rect 13245 3460 13295 3475
rect 13335 3460 13385 3475
rect 13425 3460 13475 3475
rect 13515 3460 13565 3475
rect 13605 3460 13655 3475
rect 13695 3460 13745 3475
rect 13785 3460 13835 3475
rect 13875 3460 13925 3475
rect 13965 3460 14015 3475
rect 14055 3460 14105 3475
rect 14145 3460 14195 3475
rect 14235 3460 14285 3475
rect 14325 3460 14375 3475
rect 14415 3460 14465 3475
rect 14505 3460 14555 3475
rect 14595 3460 14645 3475
rect 14685 3460 14735 3475
rect 14775 3460 14825 3475
rect 14865 3460 14915 3475
rect 14955 3460 15005 3475
rect 15045 3460 15095 3475
rect 15135 3460 15185 3475
rect 15225 3460 15275 3475
rect 15315 3460 15365 3475
rect 15405 3460 15455 3475
rect 15495 3460 15545 3475
rect 15585 3460 15635 3475
rect 15675 3460 15725 3475
rect 15765 3460 15815 3475
rect 15855 3460 15905 3475
rect 15945 3460 15995 3475
rect 16035 3460 16085 3475
rect 16125 3460 16175 3475
rect 16215 3460 16265 3475
rect 16305 3460 16355 3475
rect 16395 3460 16445 3475
rect 16485 3460 16535 3475
rect 16575 3460 16625 3475
rect 16665 3460 16715 3475
rect 16755 3460 16805 3475
rect 16845 3460 16895 3475
rect 16935 3460 16985 3475
rect 17025 3460 17075 3475
rect 17115 3460 17165 3475
rect 17205 3460 17255 3475
rect 17295 3460 17345 3475
rect 17385 3460 17435 3475
rect 17475 3460 17525 3475
rect 17565 3460 17615 3475
rect 17655 3460 17705 3475
rect 17745 3460 17795 3475
rect 17835 3460 17885 3475
rect 17925 3460 17975 3475
rect 18015 3460 18065 3475
rect 18105 3460 18155 3475
rect 18195 3460 18245 3475
rect 18285 3460 18335 3475
rect 18375 3460 18425 3475
rect 18465 3460 18515 3475
rect 18555 3460 18605 3475
rect 18645 3460 18695 3475
rect 18735 3460 18785 3475
rect 18825 3460 18875 3475
rect 18915 3460 18965 3475
rect 19005 3460 19055 3475
rect 19095 3460 19145 3475
rect 19185 3460 19235 3475
rect 19275 3460 19325 3475
rect 19365 3460 19415 3475
rect 19455 3460 19505 3475
rect 19545 3460 19595 3475
rect 19635 3460 19685 3475
rect 19725 3460 19775 3475
rect 19815 3460 19865 3475
rect 19905 3460 19955 3475
rect 19995 3460 20045 3475
rect 20085 3460 20135 3475
rect 20175 3460 20225 3475
rect 20265 3460 20315 3475
rect 20355 3460 20405 3475
rect 20445 3460 20495 3475
rect 20535 3460 20585 3475
rect 20625 3460 20675 3475
<< polycont >>
rect 9210 4170 9230 4190
rect 9300 4170 9320 4190
rect 9390 4170 9410 4190
rect 9480 4170 9500 4190
rect 9570 4170 9590 4190
rect 9660 4170 9680 4190
rect 9750 4170 9770 4190
rect 9840 4170 9860 4190
rect 9930 4170 9950 4190
rect 10020 4170 10040 4190
rect 10110 4170 10130 4190
rect 10200 4170 10220 4190
rect 10290 4170 10310 4190
rect 10380 4170 10400 4190
rect 10470 4170 10490 4190
rect 10560 4170 10580 4190
rect 10650 4170 10670 4190
rect 10740 4170 10760 4190
rect 10830 4170 10850 4190
rect 10920 4170 10940 4190
rect 11010 4170 11030 4190
rect 11100 4170 11120 4190
rect 11190 4170 11210 4190
rect 11280 4170 11300 4190
rect 11370 4170 11390 4190
rect 11460 4170 11480 4190
rect 11550 4170 11570 4190
rect 11640 4170 11660 4190
rect 11730 4170 11750 4190
rect 11820 4170 11840 4190
rect 11910 4170 11930 4190
rect 12000 4170 12020 4190
rect 12090 4170 12110 4190
rect 12180 4170 12200 4190
rect 12270 4170 12290 4190
rect 12360 4170 12380 4190
rect 12450 4170 12470 4190
rect 12540 4170 12560 4190
rect 12630 4170 12650 4190
rect 12720 4170 12740 4190
rect 12810 4170 12830 4190
rect 12900 4170 12920 4190
rect 12990 4170 13010 4190
rect 13080 4170 13100 4190
rect 13170 4170 13190 4190
rect 13260 4170 13280 4190
rect 13350 4170 13370 4190
rect 13440 4170 13460 4190
rect 13530 4170 13550 4190
rect 13620 4170 13640 4190
rect 13710 4170 13730 4190
rect 13800 4170 13820 4190
rect 13890 4170 13910 4190
rect 13980 4170 14000 4190
rect 14070 4170 14090 4190
rect 14160 4170 14180 4190
rect 14250 4170 14270 4190
rect 14340 4170 14360 4190
rect 14430 4170 14450 4190
rect 14520 4170 14540 4190
rect 14610 4170 14630 4190
rect 14700 4170 14720 4190
rect 14790 4170 14810 4190
rect 14880 4170 14900 4190
rect 14970 4170 14990 4190
rect 15060 4170 15080 4190
rect 15150 4170 15170 4190
rect 15240 4170 15260 4190
rect 15330 4170 15350 4190
rect 15420 4170 15440 4190
rect 15510 4170 15530 4190
rect 15600 4170 15620 4190
rect 15690 4170 15710 4190
rect 15780 4170 15800 4190
rect 15870 4170 15890 4190
rect 15960 4170 15980 4190
rect 16050 4170 16070 4190
rect 16140 4170 16160 4190
rect 16230 4170 16250 4190
rect 16320 4170 16340 4190
rect 16410 4170 16430 4190
rect 16500 4170 16520 4190
rect 16590 4170 16610 4190
rect 16680 4170 16700 4190
rect 16770 4170 16790 4190
rect 16860 4170 16880 4190
rect 16950 4170 16970 4190
rect 17040 4170 17060 4190
rect 17130 4170 17150 4190
rect 17220 4170 17240 4190
rect 17310 4170 17330 4190
rect 17400 4170 17420 4190
rect 17490 4170 17510 4190
rect 17580 4170 17600 4190
rect 17670 4170 17690 4190
rect 17760 4170 17780 4190
rect 17850 4170 17870 4190
rect 17940 4170 17960 4190
rect 18030 4170 18050 4190
rect 18120 4170 18140 4190
rect 18210 4170 18230 4190
rect 18300 4170 18320 4190
rect 18390 4170 18410 4190
rect 18480 4170 18500 4190
rect 18570 4170 18590 4190
rect 18660 4170 18680 4190
rect 18750 4170 18770 4190
rect 18840 4170 18860 4190
rect 18930 4170 18950 4190
rect 19020 4170 19040 4190
rect 19110 4170 19130 4190
rect 19200 4170 19220 4190
rect 19290 4170 19310 4190
rect 19380 4170 19400 4190
rect 19470 4170 19490 4190
rect 19560 4170 19580 4190
rect 19650 4170 19670 4190
rect 19740 4170 19760 4190
rect 19830 4170 19850 4190
rect 19920 4170 19940 4190
rect 20010 4170 20030 4190
rect 20100 4170 20120 4190
rect 20190 4170 20210 4190
rect 20280 4170 20300 4190
rect 20370 4170 20390 4190
rect 20460 4170 20480 4190
rect 20550 4170 20570 4190
rect 20640 4170 20660 4190
rect 9210 3600 9230 3620
rect 9300 3600 9320 3620
rect 9390 3600 9410 3620
rect 9480 3600 9500 3620
rect 9570 3600 9590 3620
rect 9660 3600 9680 3620
rect 9750 3600 9770 3620
rect 9840 3600 9860 3620
rect 9930 3600 9950 3620
rect 10020 3600 10040 3620
rect 10110 3600 10130 3620
rect 10200 3600 10220 3620
rect 10290 3600 10310 3620
rect 10380 3600 10400 3620
rect 10470 3600 10490 3620
rect 10560 3600 10580 3620
rect 10650 3600 10670 3620
rect 10740 3600 10760 3620
rect 10830 3600 10850 3620
rect 10920 3600 10940 3620
rect 11010 3600 11030 3620
rect 11100 3600 11120 3620
rect 11190 3600 11210 3620
rect 11280 3600 11300 3620
rect 11370 3600 11390 3620
rect 11460 3600 11480 3620
rect 11550 3600 11570 3620
rect 11640 3600 11660 3620
rect 11730 3600 11750 3620
rect 11820 3600 11840 3620
rect 11910 3600 11930 3620
rect 12000 3600 12020 3620
rect 12090 3600 12110 3620
rect 12180 3600 12200 3620
rect 12270 3600 12290 3620
rect 12360 3600 12380 3620
rect 12450 3600 12470 3620
rect 12540 3600 12560 3620
rect 12630 3600 12650 3620
rect 12720 3600 12740 3620
rect 12810 3600 12830 3620
rect 12900 3600 12920 3620
rect 12990 3600 13010 3620
rect 13080 3600 13100 3620
rect 13170 3600 13190 3620
rect 13260 3600 13280 3620
rect 13350 3600 13370 3620
rect 13440 3600 13460 3620
rect 13530 3600 13550 3620
rect 13620 3600 13640 3620
rect 13710 3600 13730 3620
rect 13800 3600 13820 3620
rect 13890 3600 13910 3620
rect 13980 3600 14000 3620
rect 14070 3600 14090 3620
rect 14160 3600 14180 3620
rect 14250 3600 14270 3620
rect 14340 3600 14360 3620
rect 14430 3600 14450 3620
rect 14520 3600 14540 3620
rect 14610 3600 14630 3620
rect 14700 3600 14720 3620
rect 14790 3600 14810 3620
rect 14880 3600 14900 3620
rect 14970 3600 14990 3620
rect 15060 3600 15080 3620
rect 15150 3600 15170 3620
rect 15240 3600 15260 3620
rect 15330 3600 15350 3620
rect 15420 3600 15440 3620
rect 15510 3600 15530 3620
rect 15600 3600 15620 3620
rect 15690 3600 15710 3620
rect 15780 3600 15800 3620
rect 15870 3600 15890 3620
rect 15960 3600 15980 3620
rect 16050 3600 16070 3620
rect 16140 3600 16160 3620
rect 16230 3600 16250 3620
rect 16320 3600 16340 3620
rect 16410 3600 16430 3620
rect 16500 3600 16520 3620
rect 16590 3600 16610 3620
rect 16680 3600 16700 3620
rect 16770 3600 16790 3620
rect 16860 3600 16880 3620
rect 16950 3600 16970 3620
rect 17040 3600 17060 3620
rect 17130 3600 17150 3620
rect 17220 3600 17240 3620
rect 17310 3600 17330 3620
rect 17400 3600 17420 3620
rect 17490 3600 17510 3620
rect 17580 3600 17600 3620
rect 17670 3600 17690 3620
rect 17760 3600 17780 3620
rect 17850 3600 17870 3620
rect 17940 3600 17960 3620
rect 18030 3600 18050 3620
rect 18120 3600 18140 3620
rect 18210 3600 18230 3620
rect 18300 3600 18320 3620
rect 18390 3600 18410 3620
rect 18480 3600 18500 3620
rect 18570 3600 18590 3620
rect 18660 3600 18680 3620
rect 18750 3600 18770 3620
rect 18840 3600 18860 3620
rect 18930 3600 18950 3620
rect 19020 3600 19040 3620
rect 19110 3600 19130 3620
rect 19200 3600 19220 3620
rect 19290 3600 19310 3620
rect 19380 3600 19400 3620
rect 19470 3600 19490 3620
rect 19560 3600 19580 3620
rect 19650 3600 19670 3620
rect 19740 3600 19760 3620
rect 19830 3600 19850 3620
rect 19920 3600 19940 3620
rect 20010 3600 20030 3620
rect 20100 3600 20120 3620
rect 20190 3600 20210 3620
rect 20280 3600 20300 3620
rect 20370 3600 20390 3620
rect 20460 3600 20480 3620
rect 20550 3600 20570 3620
rect 20640 3600 20660 3620
<< locali >>
rect 9030 4065 9050 4375
rect 9105 4345 9165 4365
rect 9185 4345 9210 4365
rect 9230 4345 9300 4365
rect 9320 4345 9390 4365
rect 9410 4345 9480 4365
rect 9500 4345 9570 4365
rect 9590 4345 9660 4365
rect 9680 4345 9750 4365
rect 9770 4345 9840 4365
rect 9860 4345 9885 4365
rect 9905 4345 9930 4365
rect 9950 4345 10020 4365
rect 10040 4345 10065 4365
rect 10085 4345 10110 4365
rect 10130 4345 10200 4365
rect 10220 4345 10245 4365
rect 10265 4345 10290 4365
rect 10310 4345 10380 4365
rect 10400 4345 10425 4365
rect 10445 4345 10470 4365
rect 10490 4345 10560 4365
rect 10580 4345 10605 4365
rect 10625 4345 10650 4365
rect 10670 4345 10740 4365
rect 10760 4345 10785 4365
rect 10805 4345 10830 4365
rect 10850 4345 10920 4365
rect 10940 4345 10965 4365
rect 10985 4345 11010 4365
rect 11030 4345 11100 4365
rect 11120 4345 11145 4365
rect 11165 4345 11190 4365
rect 11210 4345 11280 4365
rect 11300 4345 11325 4365
rect 11345 4345 11370 4365
rect 11390 4345 11460 4365
rect 11480 4345 11505 4365
rect 11525 4345 11550 4365
rect 11570 4345 11640 4365
rect 11660 4345 11685 4365
rect 11705 4345 11730 4365
rect 11750 4345 11820 4365
rect 11840 4345 11865 4365
rect 11885 4345 11910 4365
rect 11930 4345 12000 4365
rect 12020 4345 12045 4365
rect 12065 4345 12090 4365
rect 12110 4345 12180 4365
rect 12200 4345 12225 4365
rect 12245 4345 12270 4365
rect 12290 4345 12360 4365
rect 12380 4345 12405 4365
rect 12425 4345 12450 4365
rect 12470 4345 12540 4365
rect 12560 4345 12585 4365
rect 12605 4345 12630 4365
rect 12650 4345 12720 4365
rect 12740 4345 12765 4365
rect 12785 4345 12810 4365
rect 12830 4345 12900 4365
rect 12920 4345 12945 4365
rect 12965 4345 12990 4365
rect 13010 4345 13080 4365
rect 13100 4345 13125 4365
rect 13145 4345 13170 4365
rect 13190 4345 13260 4365
rect 13280 4345 13305 4365
rect 13325 4345 13350 4365
rect 13370 4345 13440 4365
rect 13460 4345 13485 4365
rect 13505 4345 13530 4365
rect 13550 4345 13620 4365
rect 13640 4345 13665 4365
rect 13685 4345 13710 4365
rect 13730 4345 13800 4365
rect 13820 4345 13845 4365
rect 13865 4345 13890 4365
rect 13910 4345 13980 4365
rect 14000 4345 14025 4365
rect 14045 4345 14070 4365
rect 14090 4345 14160 4365
rect 14180 4345 14205 4365
rect 14225 4345 14250 4365
rect 14270 4345 14340 4365
rect 14360 4345 14385 4365
rect 14405 4345 14430 4365
rect 14450 4345 14520 4365
rect 14540 4345 14565 4365
rect 14585 4345 14610 4365
rect 14630 4345 14700 4365
rect 14720 4345 14745 4365
rect 14765 4345 14790 4365
rect 14810 4345 14880 4365
rect 14900 4345 14925 4365
rect 14945 4345 14970 4365
rect 14990 4345 15060 4365
rect 15080 4345 15105 4365
rect 15125 4345 15150 4365
rect 15170 4345 15240 4365
rect 15260 4345 15285 4365
rect 15305 4345 15330 4365
rect 15350 4345 15420 4365
rect 15440 4345 15465 4365
rect 15485 4345 15510 4365
rect 15530 4345 15600 4365
rect 15620 4345 15645 4365
rect 15665 4345 15690 4365
rect 15710 4345 15780 4365
rect 15800 4345 15825 4365
rect 15845 4345 15870 4365
rect 15890 4345 15960 4365
rect 15980 4345 16005 4365
rect 16025 4345 16050 4365
rect 16070 4345 16140 4365
rect 16160 4345 16185 4365
rect 16205 4345 16230 4365
rect 16250 4345 16320 4365
rect 16340 4345 16365 4365
rect 16385 4345 16410 4365
rect 16430 4345 16500 4365
rect 16520 4345 16545 4365
rect 16565 4345 16590 4365
rect 16610 4345 16680 4365
rect 16700 4345 16725 4365
rect 16745 4345 16770 4365
rect 16790 4345 16860 4365
rect 16880 4345 16905 4365
rect 16925 4345 16950 4365
rect 16970 4345 17040 4365
rect 17060 4345 17085 4365
rect 17105 4345 17130 4365
rect 17150 4345 17220 4365
rect 17240 4345 17265 4365
rect 17285 4345 17310 4365
rect 17330 4345 17400 4365
rect 17420 4345 17445 4365
rect 17465 4345 17490 4365
rect 17510 4345 17580 4365
rect 17600 4345 17625 4365
rect 17645 4345 17670 4365
rect 17690 4345 17760 4365
rect 17780 4345 17805 4365
rect 17825 4345 17850 4365
rect 17870 4345 17940 4365
rect 17960 4345 17985 4365
rect 18005 4345 18030 4365
rect 18050 4345 18120 4365
rect 18140 4345 18165 4365
rect 18185 4345 18210 4365
rect 18230 4345 18300 4365
rect 18320 4345 18345 4365
rect 18365 4345 18390 4365
rect 18410 4345 18480 4365
rect 18500 4345 18525 4365
rect 18545 4345 18570 4365
rect 18590 4345 18660 4365
rect 18680 4345 18705 4365
rect 18725 4345 18750 4365
rect 18770 4345 18840 4365
rect 18860 4345 18885 4365
rect 18905 4345 18930 4365
rect 18950 4345 19020 4365
rect 19040 4345 19065 4365
rect 19085 4345 19110 4365
rect 19130 4345 19200 4365
rect 19220 4345 19245 4365
rect 19265 4345 19290 4365
rect 19310 4345 19380 4365
rect 19400 4345 19425 4365
rect 19445 4345 19470 4365
rect 19490 4345 19560 4365
rect 19580 4345 19605 4365
rect 19625 4345 19650 4365
rect 19670 4345 19740 4365
rect 19760 4345 19785 4365
rect 19805 4345 19830 4365
rect 19850 4345 19920 4365
rect 19940 4345 19965 4365
rect 19985 4345 20010 4365
rect 20030 4345 20100 4365
rect 20120 4345 20190 4365
rect 20210 4345 20280 4365
rect 20300 4345 20370 4365
rect 20390 4345 20460 4365
rect 20480 4345 20550 4365
rect 20570 4345 20640 4365
rect 20660 4345 20685 4365
rect 20705 4345 20765 4365
rect 9105 4145 9125 4345
rect 9165 4305 9185 4315
rect 9165 4215 9185 4225
rect 9255 4305 9275 4315
rect 9255 4215 9275 4225
rect 9345 4305 9365 4315
rect 9345 4215 9365 4225
rect 9435 4305 9455 4315
rect 9435 4190 9455 4225
rect 9525 4305 9545 4315
rect 9525 4215 9545 4225
rect 9615 4305 9635 4315
rect 9615 4190 9635 4225
rect 9705 4305 9725 4315
rect 9705 4215 9725 4225
rect 9795 4305 9815 4315
rect 9795 4215 9815 4225
rect 9885 4305 9905 4315
rect 9885 4215 9905 4225
rect 9975 4305 9995 4315
rect 9975 4215 9995 4225
rect 10065 4305 10085 4315
rect 10065 4215 10085 4225
rect 10155 4305 10175 4315
rect 10155 4215 10175 4225
rect 10245 4305 10265 4315
rect 10245 4215 10265 4225
rect 10335 4305 10355 4315
rect 10335 4215 10355 4225
rect 10425 4305 10445 4315
rect 10425 4215 10445 4225
rect 10515 4305 10535 4315
rect 10515 4215 10535 4225
rect 10605 4305 10625 4315
rect 10605 4215 10625 4225
rect 10695 4305 10715 4315
rect 10695 4215 10715 4225
rect 10785 4305 10805 4315
rect 10785 4215 10805 4225
rect 10875 4305 10895 4315
rect 10875 4215 10895 4225
rect 10965 4305 10985 4315
rect 10965 4215 10985 4225
rect 11055 4305 11075 4315
rect 11055 4215 11075 4225
rect 11145 4305 11165 4315
rect 11145 4215 11165 4225
rect 11235 4305 11255 4315
rect 11235 4215 11255 4225
rect 11325 4305 11345 4315
rect 11325 4215 11345 4225
rect 11415 4305 11435 4315
rect 11415 4215 11435 4225
rect 11505 4305 11525 4315
rect 11505 4215 11525 4225
rect 11595 4305 11615 4315
rect 11595 4215 11615 4225
rect 11685 4305 11705 4315
rect 11685 4215 11705 4225
rect 11775 4305 11795 4315
rect 11775 4215 11795 4225
rect 11865 4305 11885 4315
rect 11865 4215 11885 4225
rect 11955 4305 11975 4315
rect 11955 4215 11975 4225
rect 12045 4305 12065 4315
rect 12045 4215 12065 4225
rect 12135 4305 12155 4315
rect 12135 4215 12155 4225
rect 12225 4305 12245 4315
rect 12225 4215 12245 4225
rect 12315 4305 12335 4315
rect 12315 4215 12335 4225
rect 12405 4305 12425 4315
rect 12405 4215 12425 4225
rect 12495 4305 12515 4315
rect 12495 4215 12515 4225
rect 12585 4305 12605 4315
rect 12585 4215 12605 4225
rect 12675 4305 12695 4315
rect 12675 4215 12695 4225
rect 12765 4305 12785 4315
rect 12765 4215 12785 4225
rect 12855 4305 12875 4315
rect 12855 4215 12875 4225
rect 12945 4305 12965 4315
rect 12945 4215 12965 4225
rect 13035 4305 13055 4315
rect 13035 4215 13055 4225
rect 13125 4305 13145 4315
rect 13125 4215 13145 4225
rect 13215 4305 13235 4315
rect 13215 4215 13235 4225
rect 13305 4305 13325 4315
rect 13305 4215 13325 4225
rect 13395 4305 13415 4315
rect 13395 4215 13415 4225
rect 13485 4305 13505 4315
rect 13485 4215 13505 4225
rect 13575 4305 13595 4315
rect 13575 4215 13595 4225
rect 13665 4305 13685 4315
rect 13665 4215 13685 4225
rect 13755 4305 13775 4315
rect 13755 4215 13775 4225
rect 13845 4305 13865 4315
rect 13845 4215 13865 4225
rect 13935 4305 13955 4315
rect 13935 4215 13955 4225
rect 14025 4305 14045 4315
rect 14025 4215 14045 4225
rect 14115 4305 14135 4315
rect 14115 4215 14135 4225
rect 14205 4305 14225 4315
rect 14205 4215 14225 4225
rect 14295 4305 14315 4315
rect 14295 4215 14315 4225
rect 14385 4305 14405 4315
rect 14385 4215 14405 4225
rect 14475 4305 14495 4315
rect 14475 4215 14495 4225
rect 14565 4305 14585 4315
rect 14565 4215 14585 4225
rect 14655 4305 14675 4315
rect 14655 4215 14675 4225
rect 14745 4305 14765 4315
rect 14745 4215 14765 4225
rect 14835 4305 14855 4315
rect 14835 4215 14855 4225
rect 14925 4305 14945 4315
rect 14925 4215 14945 4225
rect 15015 4305 15035 4315
rect 15015 4215 15035 4225
rect 15105 4305 15125 4315
rect 15105 4215 15125 4225
rect 15195 4305 15215 4315
rect 15195 4215 15215 4225
rect 15285 4305 15305 4315
rect 15285 4215 15305 4225
rect 15375 4305 15395 4315
rect 15375 4215 15395 4225
rect 15465 4305 15485 4315
rect 15465 4215 15485 4225
rect 15555 4305 15575 4315
rect 15555 4215 15575 4225
rect 15645 4305 15665 4315
rect 15645 4215 15665 4225
rect 15735 4305 15755 4315
rect 15735 4215 15755 4225
rect 15825 4305 15845 4315
rect 15825 4215 15845 4225
rect 15915 4305 15935 4315
rect 15915 4215 15935 4225
rect 16005 4305 16025 4315
rect 16005 4215 16025 4225
rect 16095 4305 16115 4315
rect 16095 4215 16115 4225
rect 16185 4305 16205 4315
rect 16185 4215 16205 4225
rect 16275 4305 16295 4315
rect 16275 4215 16295 4225
rect 16365 4305 16385 4315
rect 16365 4215 16385 4225
rect 16455 4305 16475 4315
rect 16455 4215 16475 4225
rect 16545 4305 16565 4315
rect 16545 4215 16565 4225
rect 16635 4305 16655 4315
rect 16635 4215 16655 4225
rect 16725 4305 16745 4315
rect 16725 4215 16745 4225
rect 16815 4305 16835 4315
rect 16815 4215 16835 4225
rect 16905 4305 16925 4315
rect 16905 4215 16925 4225
rect 16995 4305 17015 4315
rect 16995 4215 17015 4225
rect 17085 4305 17105 4315
rect 17085 4215 17105 4225
rect 17175 4305 17195 4315
rect 17175 4215 17195 4225
rect 17265 4305 17285 4315
rect 17265 4215 17285 4225
rect 17355 4305 17375 4315
rect 17355 4215 17375 4225
rect 17445 4305 17465 4315
rect 17445 4215 17465 4225
rect 17535 4305 17555 4315
rect 17535 4215 17555 4225
rect 17625 4305 17645 4315
rect 17625 4215 17645 4225
rect 17715 4305 17735 4315
rect 17715 4215 17735 4225
rect 17805 4305 17825 4315
rect 17805 4215 17825 4225
rect 17895 4305 17915 4315
rect 17895 4215 17915 4225
rect 17985 4305 18005 4315
rect 17985 4215 18005 4225
rect 18075 4305 18095 4315
rect 18075 4215 18095 4225
rect 18165 4305 18185 4315
rect 18165 4215 18185 4225
rect 18255 4305 18275 4315
rect 18255 4215 18275 4225
rect 18345 4305 18365 4315
rect 18345 4215 18365 4225
rect 18435 4305 18455 4315
rect 18435 4215 18455 4225
rect 18525 4305 18545 4315
rect 18525 4215 18545 4225
rect 18615 4305 18635 4315
rect 18615 4215 18635 4225
rect 18705 4305 18725 4315
rect 18705 4215 18725 4225
rect 18795 4305 18815 4315
rect 18795 4215 18815 4225
rect 18885 4305 18905 4315
rect 18885 4215 18905 4225
rect 18975 4305 18995 4315
rect 18975 4215 18995 4225
rect 19065 4305 19085 4315
rect 19065 4215 19085 4225
rect 19155 4305 19175 4315
rect 19155 4215 19175 4225
rect 19245 4305 19265 4315
rect 19245 4215 19265 4225
rect 19335 4305 19355 4315
rect 19335 4215 19355 4225
rect 19425 4305 19445 4315
rect 19425 4215 19445 4225
rect 19515 4305 19535 4315
rect 19515 4215 19535 4225
rect 19605 4305 19625 4315
rect 19605 4215 19625 4225
rect 19695 4305 19715 4315
rect 19695 4215 19715 4225
rect 19785 4305 19805 4315
rect 19785 4215 19805 4225
rect 19875 4305 19895 4315
rect 19875 4215 19895 4225
rect 19965 4305 19985 4315
rect 19965 4215 19985 4225
rect 20055 4305 20075 4315
rect 20055 4215 20075 4225
rect 20145 4305 20165 4315
rect 20145 4215 20165 4225
rect 20235 4305 20255 4315
rect 20235 4190 20255 4225
rect 20325 4305 20345 4315
rect 20325 4215 20345 4225
rect 20415 4305 20435 4315
rect 20415 4190 20435 4225
rect 20505 4305 20525 4315
rect 20505 4215 20525 4225
rect 20595 4305 20615 4315
rect 20595 4215 20615 4225
rect 20685 4305 20705 4315
rect 20685 4215 20705 4225
rect 9200 4170 9210 4190
rect 9230 4170 9300 4190
rect 9320 4170 9390 4190
rect 9410 4170 9480 4190
rect 9500 4170 9570 4190
rect 9590 4170 9660 4190
rect 9680 4170 9750 4190
rect 9770 4170 9840 4190
rect 9860 4170 9875 4190
rect 9920 4170 9930 4190
rect 9950 4170 10020 4190
rect 10040 4170 10050 4190
rect 10100 4170 10110 4190
rect 10130 4170 10200 4190
rect 10220 4170 10230 4190
rect 10280 4170 10290 4190
rect 10310 4170 10380 4190
rect 10400 4170 10410 4190
rect 10460 4170 10470 4190
rect 10490 4170 10560 4190
rect 10580 4170 10590 4190
rect 10640 4170 10650 4190
rect 10670 4170 10740 4190
rect 10760 4170 10770 4190
rect 10820 4170 10830 4190
rect 10850 4170 10920 4190
rect 10940 4170 10950 4190
rect 11000 4170 11010 4190
rect 11030 4170 11100 4190
rect 11120 4170 11130 4190
rect 11180 4170 11190 4190
rect 11210 4170 11280 4190
rect 11300 4170 11310 4190
rect 11360 4170 11370 4190
rect 11390 4170 11460 4190
rect 11480 4170 11490 4190
rect 11540 4170 11550 4190
rect 11570 4170 11640 4190
rect 11660 4170 11670 4190
rect 11720 4170 11730 4190
rect 11750 4170 11820 4190
rect 11840 4170 11850 4190
rect 11900 4170 11910 4190
rect 11930 4170 12000 4190
rect 12020 4170 12030 4190
rect 12080 4170 12090 4190
rect 12110 4170 12180 4190
rect 12200 4170 12210 4190
rect 12260 4170 12270 4190
rect 12290 4170 12360 4190
rect 12380 4170 12390 4190
rect 12440 4170 12450 4190
rect 12470 4170 12540 4190
rect 12560 4170 12570 4190
rect 12620 4170 12630 4190
rect 12650 4170 12720 4190
rect 12740 4170 12750 4190
rect 12800 4170 12810 4190
rect 12830 4170 12900 4190
rect 12920 4170 12930 4190
rect 12980 4170 12990 4190
rect 13010 4170 13080 4190
rect 13100 4170 13110 4190
rect 13160 4170 13170 4190
rect 13190 4170 13260 4190
rect 13280 4170 13290 4190
rect 13340 4170 13350 4190
rect 13370 4170 13440 4190
rect 13460 4170 13470 4190
rect 13520 4170 13530 4190
rect 13550 4170 13620 4190
rect 13640 4170 13650 4190
rect 13700 4170 13710 4190
rect 13730 4170 13800 4190
rect 13820 4170 13830 4190
rect 13880 4170 13890 4190
rect 13910 4170 13980 4190
rect 14000 4170 14010 4190
rect 14060 4170 14070 4190
rect 14090 4170 14160 4190
rect 14180 4170 14190 4190
rect 14240 4170 14250 4190
rect 14270 4170 14340 4190
rect 14360 4170 14370 4190
rect 14420 4170 14430 4190
rect 14450 4170 14520 4190
rect 14540 4170 14550 4190
rect 14600 4170 14610 4190
rect 14630 4170 14700 4190
rect 14720 4170 14730 4190
rect 14780 4170 14790 4190
rect 14810 4170 14880 4190
rect 14900 4170 14910 4190
rect 14960 4170 14970 4190
rect 14990 4170 15060 4190
rect 15080 4170 15090 4190
rect 15140 4170 15150 4190
rect 15170 4170 15240 4190
rect 15260 4170 15270 4190
rect 15320 4170 15330 4190
rect 15350 4170 15420 4190
rect 15440 4170 15450 4190
rect 15500 4170 15510 4190
rect 15530 4170 15600 4190
rect 15620 4170 15630 4190
rect 15680 4170 15690 4190
rect 15710 4170 15780 4190
rect 15800 4170 15810 4190
rect 15860 4170 15870 4190
rect 15890 4170 15960 4190
rect 15980 4170 15990 4190
rect 16040 4170 16050 4190
rect 16070 4170 16140 4190
rect 16160 4170 16170 4190
rect 16220 4170 16230 4190
rect 16250 4170 16320 4190
rect 16340 4170 16350 4190
rect 16400 4170 16410 4190
rect 16430 4170 16500 4190
rect 16520 4170 16530 4190
rect 16580 4170 16590 4190
rect 16610 4170 16680 4190
rect 16700 4170 16710 4190
rect 16760 4170 16770 4190
rect 16790 4170 16860 4190
rect 16880 4170 16890 4190
rect 16940 4170 16950 4190
rect 16970 4170 17040 4190
rect 17060 4170 17070 4190
rect 17120 4170 17130 4190
rect 17150 4170 17220 4190
rect 17240 4170 17250 4190
rect 17300 4170 17310 4190
rect 17330 4170 17400 4190
rect 17420 4170 17430 4190
rect 17480 4170 17490 4190
rect 17510 4170 17580 4190
rect 17600 4170 17610 4190
rect 17660 4170 17670 4190
rect 17690 4170 17760 4190
rect 17780 4170 17790 4190
rect 17840 4170 17850 4190
rect 17870 4170 17940 4190
rect 17960 4170 17970 4190
rect 18020 4170 18030 4190
rect 18050 4170 18120 4190
rect 18140 4170 18150 4190
rect 18200 4170 18210 4190
rect 18230 4170 18300 4190
rect 18320 4170 18330 4190
rect 18380 4170 18390 4190
rect 18410 4170 18480 4190
rect 18500 4170 18510 4190
rect 18560 4170 18570 4190
rect 18590 4170 18660 4190
rect 18680 4170 18690 4190
rect 18740 4170 18750 4190
rect 18770 4170 18840 4190
rect 18860 4170 18870 4190
rect 18920 4170 18930 4190
rect 18950 4170 19020 4190
rect 19040 4170 19050 4190
rect 19100 4170 19110 4190
rect 19130 4170 19200 4190
rect 19220 4170 19230 4190
rect 19280 4170 19290 4190
rect 19310 4170 19380 4190
rect 19400 4170 19410 4190
rect 19460 4170 19470 4190
rect 19490 4170 19560 4190
rect 19580 4170 19590 4190
rect 19640 4170 19650 4190
rect 19670 4170 19740 4190
rect 19760 4170 19770 4190
rect 19820 4170 19830 4190
rect 19850 4170 19920 4190
rect 19940 4170 19950 4190
rect 19995 4170 20010 4190
rect 20030 4170 20100 4190
rect 20120 4170 20190 4190
rect 20210 4170 20280 4190
rect 20300 4170 20370 4190
rect 20390 4170 20460 4190
rect 20480 4170 20550 4190
rect 20570 4170 20640 4190
rect 20660 4170 20670 4190
rect 20745 4145 20765 4345
rect 9105 4125 9210 4145
rect 9230 4125 9300 4145
rect 9320 4125 9390 4145
rect 9410 4125 9480 4145
rect 9500 4125 9570 4145
rect 9590 4125 9660 4145
rect 9680 4125 9750 4145
rect 9770 4125 9840 4145
rect 9860 4125 9930 4145
rect 9950 4125 10020 4145
rect 10040 4125 10110 4145
rect 10130 4125 10200 4145
rect 10220 4125 10290 4145
rect 10310 4125 10380 4145
rect 10400 4125 10470 4145
rect 10490 4125 10560 4145
rect 10580 4125 10650 4145
rect 10670 4125 10740 4145
rect 10760 4125 10830 4145
rect 10850 4125 10920 4145
rect 10940 4125 11010 4145
rect 11030 4125 11100 4145
rect 11120 4125 11190 4145
rect 11210 4125 11280 4145
rect 11300 4125 11370 4145
rect 11390 4125 11460 4145
rect 11480 4125 11550 4145
rect 11570 4125 11640 4145
rect 11660 4125 11730 4145
rect 11750 4125 11820 4145
rect 11840 4125 11910 4145
rect 11930 4125 12000 4145
rect 12020 4125 12090 4145
rect 12110 4125 12180 4145
rect 12200 4125 12270 4145
rect 12290 4125 12360 4145
rect 12380 4125 12450 4145
rect 12470 4125 12540 4145
rect 12560 4125 12630 4145
rect 12650 4125 12720 4145
rect 12740 4125 12810 4145
rect 12830 4125 12900 4145
rect 12920 4125 12990 4145
rect 13010 4125 13080 4145
rect 13100 4125 13170 4145
rect 13190 4125 13260 4145
rect 13280 4125 13350 4145
rect 13370 4125 13440 4145
rect 13460 4125 13530 4145
rect 13550 4125 13620 4145
rect 13640 4125 13710 4145
rect 13730 4125 13800 4145
rect 13820 4125 13890 4145
rect 13910 4125 13980 4145
rect 14000 4125 14070 4145
rect 14090 4125 14160 4145
rect 14180 4125 14250 4145
rect 14270 4125 14340 4145
rect 14360 4125 14430 4145
rect 14450 4125 14520 4145
rect 14540 4125 14610 4145
rect 14630 4125 14700 4145
rect 14720 4125 14790 4145
rect 14810 4125 14880 4145
rect 14900 4125 14970 4145
rect 14990 4125 15060 4145
rect 15080 4125 15150 4145
rect 15170 4125 15240 4145
rect 15260 4125 15330 4145
rect 15350 4125 15420 4145
rect 15440 4125 15510 4145
rect 15530 4125 15600 4145
rect 15620 4125 15690 4145
rect 15710 4125 15780 4145
rect 15800 4125 15870 4145
rect 15890 4125 15960 4145
rect 15980 4125 16050 4145
rect 16070 4125 16140 4145
rect 16160 4125 16230 4145
rect 16250 4125 16320 4145
rect 16340 4125 16410 4145
rect 16430 4125 16500 4145
rect 16520 4125 16590 4145
rect 16610 4125 16680 4145
rect 16700 4125 16770 4145
rect 16790 4125 16860 4145
rect 16880 4125 16950 4145
rect 16970 4125 17040 4145
rect 17060 4125 17130 4145
rect 17150 4125 17220 4145
rect 17240 4125 17310 4145
rect 17330 4125 17400 4145
rect 17420 4125 17490 4145
rect 17510 4125 17580 4145
rect 17600 4125 17670 4145
rect 17690 4125 17760 4145
rect 17780 4125 17850 4145
rect 17870 4125 17940 4145
rect 17960 4125 18030 4145
rect 18050 4125 18120 4145
rect 18140 4125 18210 4145
rect 18230 4125 18300 4145
rect 18320 4125 18390 4145
rect 18410 4125 18480 4145
rect 18500 4125 18570 4145
rect 18590 4125 18660 4145
rect 18680 4125 18750 4145
rect 18770 4125 18840 4145
rect 18860 4125 18930 4145
rect 18950 4125 19020 4145
rect 19040 4125 19110 4145
rect 19130 4125 19200 4145
rect 19220 4125 19290 4145
rect 19310 4125 19380 4145
rect 19400 4125 19470 4145
rect 19490 4125 19560 4145
rect 19580 4125 19650 4145
rect 19670 4125 19740 4145
rect 19760 4125 19830 4145
rect 19850 4125 19920 4145
rect 19940 4125 20010 4145
rect 20030 4125 20100 4145
rect 20120 4125 20190 4145
rect 20210 4125 20280 4145
rect 20300 4125 20370 4145
rect 20390 4125 20460 4145
rect 20480 4125 20550 4145
rect 20570 4125 20640 4145
rect 20660 4125 20765 4145
rect 9155 4085 9795 4105
rect 9815 4085 11370 4105
rect 11390 4085 11685 4105
rect 11705 4085 11910 4105
rect 11930 4085 12090 4105
rect 12110 4085 12630 4105
rect 12650 4085 20145 4105
rect 20165 4085 20715 4105
rect 20820 4065 20840 4375
rect 9030 4045 9210 4065
rect 9230 4045 9300 4065
rect 9320 4045 9390 4065
rect 9410 4045 9480 4065
rect 9500 4045 9570 4065
rect 9590 4045 9660 4065
rect 9680 4045 9750 4065
rect 9770 4045 9840 4065
rect 9860 4045 9930 4065
rect 9950 4045 10020 4065
rect 10040 4045 10110 4065
rect 10130 4045 10200 4065
rect 10220 4045 10290 4065
rect 10310 4045 10380 4065
rect 10400 4045 10470 4065
rect 10490 4045 10560 4065
rect 10580 4045 10650 4065
rect 10670 4045 10740 4065
rect 10760 4045 10830 4065
rect 10850 4045 10920 4065
rect 10940 4045 11010 4065
rect 11030 4045 11100 4065
rect 11120 4045 11190 4065
rect 11210 4045 11280 4065
rect 11300 4045 11370 4065
rect 11390 4045 11460 4065
rect 11480 4045 11550 4065
rect 11570 4045 11640 4065
rect 11660 4045 11730 4065
rect 11750 4045 11820 4065
rect 11840 4045 11910 4065
rect 11930 4045 12000 4065
rect 12020 4045 12090 4065
rect 12110 4045 12180 4065
rect 12200 4045 12270 4065
rect 12290 4045 12360 4065
rect 12380 4045 12450 4065
rect 12470 4045 12540 4065
rect 12560 4045 12630 4065
rect 12650 4045 12720 4065
rect 12740 4045 12810 4065
rect 12830 4045 12900 4065
rect 12920 4045 12990 4065
rect 13010 4045 13080 4065
rect 13100 4045 13170 4065
rect 13190 4045 13260 4065
rect 13280 4045 13350 4065
rect 13370 4045 13440 4065
rect 13460 4045 13530 4065
rect 13550 4045 13620 4065
rect 13640 4045 13710 4065
rect 13730 4045 13800 4065
rect 13820 4045 13890 4065
rect 13910 4045 13980 4065
rect 14000 4045 14070 4065
rect 14090 4045 14160 4065
rect 14180 4045 14250 4065
rect 14270 4045 14340 4065
rect 14360 4045 14430 4065
rect 14450 4045 14520 4065
rect 14540 4045 14610 4065
rect 14630 4045 14700 4065
rect 14720 4045 14790 4065
rect 14810 4045 14880 4065
rect 14900 4045 14970 4065
rect 14990 4045 15060 4065
rect 15080 4045 15150 4065
rect 15170 4045 15240 4065
rect 15260 4045 15330 4065
rect 15350 4045 15420 4065
rect 15440 4045 15510 4065
rect 15530 4045 15600 4065
rect 15620 4045 15690 4065
rect 15710 4045 15780 4065
rect 15800 4045 15870 4065
rect 15890 4045 15960 4065
rect 15980 4045 16050 4065
rect 16070 4045 16140 4065
rect 16160 4045 16230 4065
rect 16250 4045 16320 4065
rect 16340 4045 16410 4065
rect 16430 4045 16500 4065
rect 16520 4045 16590 4065
rect 16610 4045 16680 4065
rect 16700 4045 16770 4065
rect 16790 4045 16860 4065
rect 16880 4045 16950 4065
rect 16970 4045 17040 4065
rect 17060 4045 17130 4065
rect 17150 4045 17220 4065
rect 17240 4045 17310 4065
rect 17330 4045 17400 4065
rect 17420 4045 17490 4065
rect 17510 4045 17580 4065
rect 17600 4045 17670 4065
rect 17690 4045 17760 4065
rect 17780 4045 17850 4065
rect 17870 4045 17940 4065
rect 17960 4045 18030 4065
rect 18050 4045 18120 4065
rect 18140 4045 18210 4065
rect 18230 4045 18300 4065
rect 18320 4045 18390 4065
rect 18410 4045 18480 4065
rect 18500 4045 18570 4065
rect 18590 4045 18660 4065
rect 18680 4045 18750 4065
rect 18770 4045 18840 4065
rect 18860 4045 18930 4065
rect 18950 4045 19020 4065
rect 19040 4045 19110 4065
rect 19130 4045 19200 4065
rect 19220 4045 19290 4065
rect 19310 4045 19380 4065
rect 19400 4045 19470 4065
rect 19490 4045 19560 4065
rect 19580 4045 19650 4065
rect 19670 4045 19740 4065
rect 19760 4045 19830 4065
rect 19850 4045 19920 4065
rect 19940 4045 20010 4065
rect 20030 4045 20100 4065
rect 20120 4045 20190 4065
rect 20210 4045 20280 4065
rect 20300 4045 20370 4065
rect 20390 4045 20460 4065
rect 20480 4045 20550 4065
rect 20570 4045 20640 4065
rect 20660 4045 20840 4065
rect 9155 4005 11460 4025
rect 11480 4005 12000 4025
rect 12020 4005 20715 4025
rect 9155 3965 11640 3985
rect 11660 3965 11820 3985
rect 11840 3965 20325 3985
rect 20345 3965 20715 3985
rect 9155 3925 10785 3945
rect 10805 3925 11145 3945
rect 11165 3925 12225 3945
rect 12245 3925 12585 3945
rect 12605 3925 20415 3945
rect 20435 3925 20715 3945
rect 9155 3885 12270 3905
rect 12290 3885 12360 3905
rect 12380 3885 12405 3905
rect 12425 3885 12450 3905
rect 12470 3885 12540 3905
rect 12560 3885 20235 3905
rect 20255 3885 20715 3905
rect 9155 3845 10920 3865
rect 10940 3845 11100 3865
rect 11120 3845 11550 3865
rect 11570 3845 11730 3865
rect 11750 3845 20715 3865
rect 9155 3805 11505 3825
rect 11525 3805 11865 3825
rect 11885 3805 12045 3825
rect 12065 3805 20715 3825
rect 9155 3765 10740 3785
rect 10760 3765 10965 3785
rect 10985 3765 11280 3785
rect 11300 3765 12180 3785
rect 12200 3765 12720 3785
rect 12740 3765 20715 3785
rect 9155 3725 10830 3745
rect 10850 3725 11010 3745
rect 11030 3725 20505 3745
rect 20525 3725 20715 3745
rect 9155 3685 10650 3705
rect 10670 3685 11190 3705
rect 11210 3685 20595 3705
rect 20615 3685 20715 3705
rect 9030 3645 9210 3665
rect 9230 3645 9300 3665
rect 9320 3645 9390 3665
rect 9410 3645 9480 3665
rect 9500 3645 9570 3665
rect 9590 3645 9660 3665
rect 9680 3645 9750 3665
rect 9770 3645 9840 3665
rect 9860 3645 9930 3665
rect 9950 3645 10020 3665
rect 10040 3645 10110 3665
rect 10130 3645 10200 3665
rect 10220 3645 10290 3665
rect 10310 3645 10380 3665
rect 10400 3645 10470 3665
rect 10490 3645 10560 3665
rect 10580 3645 10650 3665
rect 10670 3645 10740 3665
rect 10760 3645 10830 3665
rect 10850 3645 10920 3665
rect 10940 3645 11010 3665
rect 11030 3645 11100 3665
rect 11120 3645 11190 3665
rect 11210 3645 11280 3665
rect 11300 3645 11370 3665
rect 11390 3645 11460 3665
rect 11480 3645 11550 3665
rect 11570 3645 11640 3665
rect 11660 3645 11730 3665
rect 11750 3645 11820 3665
rect 11840 3645 11910 3665
rect 11930 3645 12000 3665
rect 12020 3645 12090 3665
rect 12110 3645 12180 3665
rect 12200 3645 12270 3665
rect 12290 3645 12360 3665
rect 12380 3645 12450 3665
rect 12470 3645 12540 3665
rect 12560 3645 12630 3665
rect 12650 3645 12720 3665
rect 12740 3645 12810 3665
rect 12830 3645 12900 3665
rect 12920 3645 12990 3665
rect 13010 3645 13080 3665
rect 13100 3645 13170 3665
rect 13190 3645 13260 3665
rect 13280 3645 13350 3665
rect 13370 3645 13440 3665
rect 13460 3645 13530 3665
rect 13550 3645 13620 3665
rect 13640 3645 13710 3665
rect 13730 3645 13800 3665
rect 13820 3645 13890 3665
rect 13910 3645 13980 3665
rect 14000 3645 14070 3665
rect 14090 3645 14160 3665
rect 14180 3645 14250 3665
rect 14270 3645 14340 3665
rect 14360 3645 14430 3665
rect 14450 3645 14520 3665
rect 14540 3645 14610 3665
rect 14630 3645 14700 3665
rect 14720 3645 14790 3665
rect 14810 3645 14880 3665
rect 14900 3645 14970 3665
rect 14990 3645 15060 3665
rect 15080 3645 15150 3665
rect 15170 3645 15240 3665
rect 15260 3645 15330 3665
rect 15350 3645 15420 3665
rect 15440 3645 15510 3665
rect 15530 3645 15600 3665
rect 15620 3645 15690 3665
rect 15710 3645 15780 3665
rect 15800 3645 15870 3665
rect 15890 3645 15960 3665
rect 15980 3645 16050 3665
rect 16070 3645 16140 3665
rect 16160 3645 16230 3665
rect 16250 3645 16320 3665
rect 16340 3645 16410 3665
rect 16430 3645 16500 3665
rect 16520 3645 16590 3665
rect 16610 3645 16680 3665
rect 16700 3645 16770 3665
rect 16790 3645 16860 3665
rect 16880 3645 16950 3665
rect 16970 3645 17040 3665
rect 17060 3645 17130 3665
rect 17150 3645 17220 3665
rect 17240 3645 17310 3665
rect 17330 3645 17400 3665
rect 17420 3645 17490 3665
rect 17510 3645 17580 3665
rect 17600 3645 17670 3665
rect 17690 3645 17760 3665
rect 17780 3645 17850 3665
rect 17870 3645 17940 3665
rect 17960 3645 18030 3665
rect 18050 3645 18120 3665
rect 18140 3645 18210 3665
rect 18230 3645 18300 3665
rect 18320 3645 18390 3665
rect 18410 3645 18480 3665
rect 18500 3645 18570 3665
rect 18590 3645 18660 3665
rect 18680 3645 18750 3665
rect 18770 3645 18840 3665
rect 18860 3645 18930 3665
rect 18950 3645 19020 3665
rect 19040 3645 19110 3665
rect 19130 3645 19200 3665
rect 19220 3645 19290 3665
rect 19310 3645 19380 3665
rect 19400 3645 19470 3665
rect 19490 3645 19560 3665
rect 19580 3645 19650 3665
rect 19670 3645 19740 3665
rect 19760 3645 19830 3665
rect 19850 3645 19920 3665
rect 19940 3645 20010 3665
rect 20030 3645 20100 3665
rect 20120 3645 20190 3665
rect 20210 3645 20280 3665
rect 20300 3645 20370 3665
rect 20390 3645 20460 3665
rect 20480 3645 20550 3665
rect 20570 3645 20640 3665
rect 20660 3645 20840 3665
rect 9030 3445 9050 3645
rect 9200 3600 9210 3620
rect 9230 3600 9300 3620
rect 9320 3600 9390 3620
rect 9410 3600 9480 3620
rect 9500 3600 9570 3620
rect 9590 3600 9660 3620
rect 9680 3600 9750 3620
rect 9770 3600 9840 3620
rect 9860 3600 9870 3620
rect 9920 3600 9930 3620
rect 9950 3600 10020 3620
rect 10040 3600 10050 3620
rect 10100 3600 10110 3620
rect 10130 3600 10200 3620
rect 10220 3600 10230 3620
rect 10280 3600 10290 3620
rect 10310 3600 10380 3620
rect 10400 3600 10410 3620
rect 10460 3600 10470 3620
rect 10490 3600 10560 3620
rect 10580 3600 10590 3620
rect 10640 3600 10650 3620
rect 10670 3600 10740 3620
rect 10760 3600 10770 3620
rect 10820 3600 10830 3620
rect 10850 3600 10920 3620
rect 10940 3600 10950 3620
rect 11000 3600 11010 3620
rect 11030 3600 11100 3620
rect 11120 3600 11130 3620
rect 11180 3600 11190 3620
rect 11210 3600 11280 3620
rect 11300 3600 11310 3620
rect 11360 3600 11370 3620
rect 11390 3600 11460 3620
rect 11480 3600 11490 3620
rect 11540 3600 11550 3620
rect 11570 3600 11640 3620
rect 11660 3600 11670 3620
rect 11720 3600 11730 3620
rect 11750 3600 11820 3620
rect 11840 3600 11850 3620
rect 11900 3600 11910 3620
rect 11930 3600 12000 3620
rect 12020 3600 12030 3620
rect 12080 3600 12090 3620
rect 12110 3600 12180 3620
rect 12200 3600 12210 3620
rect 12260 3600 12270 3620
rect 12290 3600 12360 3620
rect 12380 3600 12390 3620
rect 12440 3600 12450 3620
rect 12470 3600 12540 3620
rect 12560 3600 12570 3620
rect 12620 3600 12630 3620
rect 12650 3600 12720 3620
rect 12740 3600 12750 3620
rect 12800 3600 12810 3620
rect 12830 3600 12900 3620
rect 12920 3600 12930 3620
rect 12980 3600 12990 3620
rect 13010 3600 13080 3620
rect 13100 3600 13110 3620
rect 13160 3600 13170 3620
rect 13190 3600 13260 3620
rect 13280 3600 13290 3620
rect 13340 3600 13350 3620
rect 13370 3600 13440 3620
rect 13460 3600 13470 3620
rect 13520 3600 13530 3620
rect 13550 3600 13620 3620
rect 13640 3600 13650 3620
rect 13700 3600 13710 3620
rect 13730 3600 13800 3620
rect 13820 3600 13830 3620
rect 13880 3600 13890 3620
rect 13910 3600 13980 3620
rect 14000 3600 14010 3620
rect 14060 3600 14070 3620
rect 14090 3600 14160 3620
rect 14180 3600 14190 3620
rect 14240 3600 14250 3620
rect 14270 3600 14340 3620
rect 14360 3600 14370 3620
rect 14420 3600 14430 3620
rect 14450 3600 14520 3620
rect 14540 3600 14550 3620
rect 14600 3600 14610 3620
rect 14630 3600 14700 3620
rect 14720 3600 14730 3620
rect 14780 3600 14790 3620
rect 14810 3600 14880 3620
rect 14900 3600 14910 3620
rect 14960 3600 14970 3620
rect 14990 3600 15060 3620
rect 15080 3600 15090 3620
rect 15140 3600 15150 3620
rect 15170 3600 15240 3620
rect 15260 3600 15270 3620
rect 15320 3600 15330 3620
rect 15350 3600 15420 3620
rect 15440 3600 15450 3620
rect 15500 3600 15510 3620
rect 15530 3600 15600 3620
rect 15620 3600 15630 3620
rect 15680 3600 15690 3620
rect 15710 3600 15780 3620
rect 15800 3600 15810 3620
rect 15860 3600 15870 3620
rect 15890 3600 15960 3620
rect 15980 3600 15990 3620
rect 16040 3600 16050 3620
rect 16070 3600 16140 3620
rect 16160 3600 16170 3620
rect 16220 3600 16230 3620
rect 16250 3600 16320 3620
rect 16340 3600 16350 3620
rect 16400 3600 16410 3620
rect 16430 3600 16500 3620
rect 16520 3600 16530 3620
rect 16580 3600 16590 3620
rect 16610 3600 16680 3620
rect 16700 3600 16710 3620
rect 16760 3600 16770 3620
rect 16790 3600 16860 3620
rect 16880 3600 16890 3620
rect 16940 3600 16950 3620
rect 16970 3600 17040 3620
rect 17060 3600 17070 3620
rect 17120 3600 17130 3620
rect 17150 3600 17220 3620
rect 17240 3600 17250 3620
rect 17300 3600 17310 3620
rect 17330 3600 17400 3620
rect 17420 3600 17430 3620
rect 17480 3600 17490 3620
rect 17510 3600 17580 3620
rect 17600 3600 17610 3620
rect 17660 3600 17670 3620
rect 17690 3600 17760 3620
rect 17780 3600 17790 3620
rect 17840 3600 17850 3620
rect 17870 3600 17940 3620
rect 17960 3600 17970 3620
rect 18020 3600 18030 3620
rect 18050 3600 18120 3620
rect 18140 3600 18150 3620
rect 18200 3600 18210 3620
rect 18230 3600 18300 3620
rect 18320 3600 18330 3620
rect 18380 3600 18390 3620
rect 18410 3600 18480 3620
rect 18500 3600 18510 3620
rect 18560 3600 18570 3620
rect 18590 3600 18660 3620
rect 18680 3600 18690 3620
rect 18740 3600 18750 3620
rect 18770 3600 18840 3620
rect 18860 3600 18870 3620
rect 18920 3600 18930 3620
rect 18950 3600 19020 3620
rect 19040 3600 19050 3620
rect 19100 3600 19110 3620
rect 19130 3600 19200 3620
rect 19220 3600 19230 3620
rect 19280 3600 19290 3620
rect 19310 3600 19380 3620
rect 19400 3600 19410 3620
rect 19460 3600 19470 3620
rect 19490 3600 19560 3620
rect 19580 3600 19590 3620
rect 19640 3600 19650 3620
rect 19670 3600 19740 3620
rect 19760 3600 19770 3620
rect 19820 3600 19830 3620
rect 19850 3600 19920 3620
rect 19940 3600 19950 3620
rect 20000 3600 20010 3620
rect 20030 3600 20100 3620
rect 20120 3600 20190 3620
rect 20210 3600 20280 3620
rect 20300 3600 20370 3620
rect 20390 3600 20460 3620
rect 20480 3600 20550 3620
rect 20570 3600 20640 3620
rect 20660 3600 20670 3620
rect 9165 3565 9185 3575
rect 9165 3475 9185 3485
rect 9255 3565 9275 3575
rect 9255 3475 9275 3485
rect 9345 3565 9365 3575
rect 9345 3475 9365 3485
rect 9435 3565 9455 3600
rect 9435 3475 9455 3485
rect 9525 3565 9545 3575
rect 9525 3475 9545 3485
rect 9615 3565 9635 3600
rect 9615 3475 9635 3485
rect 9705 3565 9725 3575
rect 9705 3475 9725 3485
rect 9795 3565 9815 3575
rect 9795 3475 9815 3485
rect 9885 3565 9905 3575
rect 9885 3475 9905 3485
rect 9975 3565 9995 3575
rect 9975 3475 9995 3485
rect 10065 3565 10085 3575
rect 10065 3475 10085 3485
rect 10155 3565 10175 3575
rect 10155 3475 10175 3485
rect 10245 3565 10265 3575
rect 10245 3475 10265 3485
rect 10335 3565 10355 3575
rect 10335 3475 10355 3485
rect 10425 3565 10445 3575
rect 10425 3475 10445 3485
rect 10515 3565 10535 3575
rect 10515 3475 10535 3485
rect 10605 3565 10625 3575
rect 10605 3475 10625 3485
rect 10695 3565 10715 3575
rect 10695 3475 10715 3485
rect 10785 3565 10805 3575
rect 10785 3475 10805 3485
rect 10875 3565 10895 3575
rect 10875 3475 10895 3485
rect 10965 3565 10985 3575
rect 10965 3475 10985 3485
rect 11055 3565 11075 3575
rect 11055 3475 11075 3485
rect 11145 3565 11165 3575
rect 11145 3475 11165 3485
rect 11235 3565 11255 3575
rect 11235 3475 11255 3485
rect 11325 3565 11345 3575
rect 11325 3475 11345 3485
rect 11415 3565 11435 3575
rect 11415 3475 11435 3485
rect 11505 3565 11525 3575
rect 11505 3475 11525 3485
rect 11595 3565 11615 3575
rect 11595 3475 11615 3485
rect 11685 3565 11705 3575
rect 11685 3475 11705 3485
rect 11775 3565 11795 3575
rect 11775 3475 11795 3485
rect 11865 3565 11885 3575
rect 11865 3475 11885 3485
rect 11955 3565 11975 3575
rect 11955 3475 11975 3485
rect 12045 3565 12065 3575
rect 12045 3475 12065 3485
rect 12135 3565 12155 3575
rect 12135 3475 12155 3485
rect 12225 3565 12245 3575
rect 12225 3475 12245 3485
rect 12315 3565 12335 3575
rect 12315 3475 12335 3485
rect 12405 3565 12425 3575
rect 12405 3475 12425 3485
rect 12495 3565 12515 3575
rect 12495 3475 12515 3485
rect 12585 3565 12605 3575
rect 12585 3475 12605 3485
rect 12675 3565 12695 3575
rect 12675 3475 12695 3485
rect 12765 3565 12785 3575
rect 12765 3475 12785 3485
rect 12855 3565 12875 3575
rect 12855 3475 12875 3485
rect 12945 3565 12965 3575
rect 12945 3475 12965 3485
rect 13035 3565 13055 3575
rect 13035 3475 13055 3485
rect 13125 3565 13145 3575
rect 13125 3475 13145 3485
rect 13215 3565 13235 3575
rect 13215 3475 13235 3485
rect 13305 3565 13325 3575
rect 13305 3475 13325 3485
rect 13395 3565 13415 3575
rect 13395 3475 13415 3485
rect 13485 3565 13505 3575
rect 13485 3475 13505 3485
rect 13575 3565 13595 3575
rect 13575 3475 13595 3485
rect 13665 3565 13685 3575
rect 13665 3475 13685 3485
rect 13755 3565 13775 3575
rect 13755 3475 13775 3485
rect 13845 3565 13865 3575
rect 13845 3475 13865 3485
rect 13935 3565 13955 3575
rect 13935 3475 13955 3485
rect 14025 3565 14045 3575
rect 14025 3475 14045 3485
rect 14115 3565 14135 3575
rect 14115 3475 14135 3485
rect 14205 3565 14225 3575
rect 14205 3475 14225 3485
rect 14295 3565 14315 3575
rect 14295 3475 14315 3485
rect 14385 3565 14405 3575
rect 14385 3475 14405 3485
rect 14475 3565 14495 3575
rect 14475 3475 14495 3485
rect 14565 3565 14585 3575
rect 14565 3475 14585 3485
rect 14655 3565 14675 3575
rect 14655 3475 14675 3485
rect 14745 3565 14765 3575
rect 14745 3475 14765 3485
rect 14835 3565 14855 3575
rect 14835 3475 14855 3485
rect 14925 3565 14945 3575
rect 14925 3475 14945 3485
rect 15015 3565 15035 3575
rect 15015 3475 15035 3485
rect 15105 3565 15125 3575
rect 15105 3475 15125 3485
rect 15195 3565 15215 3575
rect 15195 3475 15215 3485
rect 15285 3565 15305 3575
rect 15285 3475 15305 3485
rect 15375 3565 15395 3575
rect 15375 3475 15395 3485
rect 15465 3565 15485 3575
rect 15465 3475 15485 3485
rect 15555 3565 15575 3575
rect 15555 3475 15575 3485
rect 15645 3565 15665 3575
rect 15645 3475 15665 3485
rect 15735 3565 15755 3575
rect 15735 3475 15755 3485
rect 15825 3565 15845 3575
rect 15825 3475 15845 3485
rect 15915 3565 15935 3575
rect 15915 3475 15935 3485
rect 16005 3565 16025 3575
rect 16005 3475 16025 3485
rect 16095 3565 16115 3575
rect 16095 3475 16115 3485
rect 16185 3565 16205 3575
rect 16185 3475 16205 3485
rect 16275 3565 16295 3575
rect 16275 3475 16295 3485
rect 16365 3565 16385 3575
rect 16365 3475 16385 3485
rect 16455 3565 16475 3575
rect 16455 3475 16475 3485
rect 16545 3565 16565 3575
rect 16545 3475 16565 3485
rect 16635 3565 16655 3575
rect 16635 3475 16655 3485
rect 16725 3565 16745 3575
rect 16725 3475 16745 3485
rect 16815 3565 16835 3575
rect 16815 3475 16835 3485
rect 16905 3565 16925 3575
rect 16905 3475 16925 3485
rect 16995 3565 17015 3575
rect 16995 3475 17015 3485
rect 17085 3565 17105 3575
rect 17085 3475 17105 3485
rect 17175 3565 17195 3575
rect 17175 3475 17195 3485
rect 17265 3565 17285 3575
rect 17265 3475 17285 3485
rect 17355 3565 17375 3575
rect 17355 3475 17375 3485
rect 17445 3565 17465 3575
rect 17445 3475 17465 3485
rect 17535 3565 17555 3575
rect 17535 3475 17555 3485
rect 17625 3565 17645 3575
rect 17625 3475 17645 3485
rect 17715 3565 17735 3575
rect 17715 3475 17735 3485
rect 17805 3565 17825 3575
rect 17805 3475 17825 3485
rect 17895 3565 17915 3575
rect 17895 3475 17915 3485
rect 17985 3565 18005 3575
rect 17985 3475 18005 3485
rect 18075 3565 18095 3575
rect 18075 3475 18095 3485
rect 18165 3565 18185 3575
rect 18165 3475 18185 3485
rect 18255 3565 18275 3575
rect 18255 3475 18275 3485
rect 18345 3565 18365 3575
rect 18345 3475 18365 3485
rect 18435 3565 18455 3575
rect 18435 3475 18455 3485
rect 18525 3565 18545 3575
rect 18525 3475 18545 3485
rect 18615 3565 18635 3575
rect 18615 3475 18635 3485
rect 18705 3565 18725 3575
rect 18705 3475 18725 3485
rect 18795 3565 18815 3575
rect 18795 3475 18815 3485
rect 18885 3565 18905 3575
rect 18885 3475 18905 3485
rect 18975 3565 18995 3575
rect 18975 3475 18995 3485
rect 19065 3565 19085 3575
rect 19065 3475 19085 3485
rect 19155 3565 19175 3575
rect 19155 3475 19175 3485
rect 19245 3565 19265 3575
rect 19245 3475 19265 3485
rect 19335 3565 19355 3575
rect 19335 3475 19355 3485
rect 19425 3565 19445 3575
rect 19425 3475 19445 3485
rect 19515 3565 19535 3575
rect 19515 3475 19535 3485
rect 19605 3565 19625 3575
rect 19605 3475 19625 3485
rect 19695 3565 19715 3575
rect 19695 3475 19715 3485
rect 19785 3565 19805 3575
rect 19785 3475 19805 3485
rect 19875 3565 19895 3575
rect 19875 3475 19895 3485
rect 19965 3565 19985 3575
rect 19965 3475 19985 3485
rect 20055 3565 20075 3575
rect 20055 3475 20075 3485
rect 20145 3565 20165 3575
rect 20145 3475 20165 3485
rect 20235 3565 20255 3600
rect 20235 3475 20255 3485
rect 20325 3565 20345 3575
rect 20325 3475 20345 3485
rect 20415 3565 20435 3600
rect 20415 3475 20435 3485
rect 20505 3565 20525 3575
rect 20505 3475 20525 3485
rect 20595 3565 20615 3575
rect 20595 3475 20615 3485
rect 20685 3565 20705 3575
rect 20685 3475 20705 3485
rect 20820 3445 20840 3645
rect 9020 3425 9030 3445
rect 9050 3425 9165 3445
rect 9185 3425 9210 3445
rect 9230 3425 9300 3445
rect 9320 3425 9390 3445
rect 9410 3425 9480 3445
rect 9500 3425 9570 3445
rect 9590 3425 9660 3445
rect 9680 3425 9750 3445
rect 9770 3425 9840 3445
rect 9860 3425 9885 3445
rect 9905 3425 9930 3445
rect 9950 3425 10020 3445
rect 10040 3425 10065 3445
rect 10085 3425 10110 3445
rect 10130 3425 10200 3445
rect 10220 3425 10245 3445
rect 10265 3425 10290 3445
rect 10310 3425 10380 3445
rect 10400 3425 10425 3445
rect 10445 3425 10470 3445
rect 10490 3425 10560 3445
rect 10580 3425 10605 3445
rect 10625 3425 10650 3445
rect 10670 3425 10740 3445
rect 10760 3425 10785 3445
rect 10805 3425 10830 3445
rect 10850 3425 10920 3445
rect 10940 3425 10965 3445
rect 10985 3425 11010 3445
rect 11030 3425 11100 3445
rect 11120 3425 11145 3445
rect 11165 3425 11190 3445
rect 11210 3425 11280 3445
rect 11300 3425 11325 3445
rect 11345 3425 11370 3445
rect 11390 3425 11460 3445
rect 11480 3425 11505 3445
rect 11525 3425 11550 3445
rect 11570 3425 11640 3445
rect 11660 3425 11685 3445
rect 11705 3425 11730 3445
rect 11750 3425 11820 3445
rect 11840 3425 11865 3445
rect 11885 3425 11910 3445
rect 11930 3425 12000 3445
rect 12020 3425 12045 3445
rect 12065 3425 12090 3445
rect 12110 3425 12180 3445
rect 12200 3425 12225 3445
rect 12245 3425 12270 3445
rect 12290 3425 12360 3445
rect 12380 3425 12405 3445
rect 12425 3425 12450 3445
rect 12470 3425 12540 3445
rect 12560 3425 12585 3445
rect 12605 3425 12630 3445
rect 12650 3425 12720 3445
rect 12740 3425 12765 3445
rect 12785 3425 12810 3445
rect 12830 3425 12900 3445
rect 12920 3425 12945 3445
rect 12965 3425 12990 3445
rect 13010 3425 13080 3445
rect 13100 3425 13125 3445
rect 13145 3425 13170 3445
rect 13190 3425 13260 3445
rect 13280 3425 13305 3445
rect 13325 3425 13350 3445
rect 13370 3425 13440 3445
rect 13460 3425 13485 3445
rect 13505 3425 13530 3445
rect 13550 3425 13620 3445
rect 13640 3425 13665 3445
rect 13685 3425 13710 3445
rect 13730 3425 13800 3445
rect 13820 3425 13845 3445
rect 13865 3425 13890 3445
rect 13910 3425 13980 3445
rect 14000 3425 14025 3445
rect 14045 3425 14070 3445
rect 14090 3425 14160 3445
rect 14180 3425 14205 3445
rect 14225 3425 14250 3445
rect 14270 3425 14340 3445
rect 14360 3425 14385 3445
rect 14405 3425 14430 3445
rect 14450 3425 14520 3445
rect 14540 3425 14565 3445
rect 14585 3425 14610 3445
rect 14630 3425 14700 3445
rect 14720 3425 14745 3445
rect 14765 3425 14790 3445
rect 14810 3425 14880 3445
rect 14900 3425 14925 3445
rect 14945 3425 14970 3445
rect 14990 3425 15060 3445
rect 15080 3425 15105 3445
rect 15125 3425 15150 3445
rect 15170 3425 15240 3445
rect 15260 3425 15285 3445
rect 15305 3425 15330 3445
rect 15350 3425 15420 3445
rect 15440 3425 15465 3445
rect 15485 3425 15510 3445
rect 15530 3425 15600 3445
rect 15620 3425 15645 3445
rect 15665 3425 15690 3445
rect 15710 3425 15780 3445
rect 15800 3425 15825 3445
rect 15845 3425 15870 3445
rect 15890 3425 15960 3445
rect 15980 3425 16005 3445
rect 16025 3425 16050 3445
rect 16070 3425 16140 3445
rect 16160 3425 16185 3445
rect 16205 3425 16230 3445
rect 16250 3425 16320 3445
rect 16340 3425 16365 3445
rect 16385 3425 16410 3445
rect 16430 3425 16500 3445
rect 16520 3425 16545 3445
rect 16565 3425 16590 3445
rect 16610 3425 16680 3445
rect 16700 3425 16725 3445
rect 16745 3425 16770 3445
rect 16790 3425 16860 3445
rect 16880 3425 16905 3445
rect 16925 3425 16950 3445
rect 16970 3425 17040 3445
rect 17060 3425 17085 3445
rect 17105 3425 17130 3445
rect 17150 3425 17220 3445
rect 17240 3425 17265 3445
rect 17285 3425 17310 3445
rect 17330 3425 17400 3445
rect 17420 3425 17445 3445
rect 17465 3425 17490 3445
rect 17510 3425 17580 3445
rect 17600 3425 17625 3445
rect 17645 3425 17670 3445
rect 17690 3425 17760 3445
rect 17780 3425 17805 3445
rect 17825 3425 17850 3445
rect 17870 3425 17940 3445
rect 17960 3425 17985 3445
rect 18005 3425 18030 3445
rect 18050 3425 18120 3445
rect 18140 3425 18165 3445
rect 18185 3425 18210 3445
rect 18230 3425 18300 3445
rect 18320 3425 18345 3445
rect 18365 3425 18390 3445
rect 18410 3425 18480 3445
rect 18500 3425 18525 3445
rect 18545 3425 18570 3445
rect 18590 3425 18660 3445
rect 18680 3425 18705 3445
rect 18725 3425 18750 3445
rect 18770 3425 18840 3445
rect 18860 3425 18885 3445
rect 18905 3425 18930 3445
rect 18950 3425 19020 3445
rect 19040 3425 19065 3445
rect 19085 3425 19110 3445
rect 19130 3425 19200 3445
rect 19220 3425 19245 3445
rect 19265 3425 19290 3445
rect 19310 3425 19380 3445
rect 19400 3425 19425 3445
rect 19445 3425 19470 3445
rect 19490 3425 19560 3445
rect 19580 3425 19605 3445
rect 19625 3425 19650 3445
rect 19670 3425 19740 3445
rect 19760 3425 19785 3445
rect 19805 3425 19830 3445
rect 19850 3425 19920 3445
rect 19940 3425 19965 3445
rect 19985 3425 20010 3445
rect 20030 3425 20100 3445
rect 20120 3425 20190 3445
rect 20210 3425 20280 3445
rect 20300 3425 20370 3445
rect 20390 3425 20460 3445
rect 20480 3425 20550 3445
rect 20570 3425 20640 3445
rect 20660 3425 20685 3445
rect 20705 3425 20820 3445
rect 20840 3425 20850 3445
<< viali >>
rect 9165 4345 9185 4365
rect 9885 4345 9905 4365
rect 10065 4345 10085 4365
rect 10245 4345 10265 4365
rect 10425 4345 10445 4365
rect 10605 4345 10625 4365
rect 10785 4345 10805 4365
rect 10965 4345 10985 4365
rect 11145 4345 11165 4365
rect 11325 4345 11345 4365
rect 11505 4345 11525 4365
rect 11685 4345 11705 4365
rect 11865 4345 11885 4365
rect 12045 4345 12065 4365
rect 12225 4345 12245 4365
rect 12405 4345 12425 4365
rect 12585 4345 12605 4365
rect 12765 4345 12785 4365
rect 12945 4345 12965 4365
rect 13125 4345 13145 4365
rect 13305 4345 13325 4365
rect 13485 4345 13505 4365
rect 13665 4345 13685 4365
rect 13845 4345 13865 4365
rect 14025 4345 14045 4365
rect 14205 4345 14225 4365
rect 14385 4345 14405 4365
rect 14565 4345 14585 4365
rect 14745 4345 14765 4365
rect 14925 4345 14945 4365
rect 15105 4345 15125 4365
rect 15285 4345 15305 4365
rect 15465 4345 15485 4365
rect 15645 4345 15665 4365
rect 15825 4345 15845 4365
rect 16005 4345 16025 4365
rect 16185 4345 16205 4365
rect 16365 4345 16385 4365
rect 16545 4345 16565 4365
rect 16725 4345 16745 4365
rect 16905 4345 16925 4365
rect 17085 4345 17105 4365
rect 17265 4345 17285 4365
rect 17445 4345 17465 4365
rect 17625 4345 17645 4365
rect 17805 4345 17825 4365
rect 17985 4345 18005 4365
rect 18165 4345 18185 4365
rect 18345 4345 18365 4365
rect 18525 4345 18545 4365
rect 18705 4345 18725 4365
rect 18885 4345 18905 4365
rect 19065 4345 19085 4365
rect 19245 4345 19265 4365
rect 19425 4345 19445 4365
rect 19605 4345 19625 4365
rect 19785 4345 19805 4365
rect 19965 4345 19985 4365
rect 20685 4345 20705 4365
rect 9165 4225 9185 4305
rect 9885 4225 9905 4305
rect 9975 4225 9995 4305
rect 10065 4225 10085 4305
rect 10155 4225 10175 4305
rect 10245 4225 10265 4305
rect 10335 4225 10355 4305
rect 10425 4225 10445 4305
rect 10515 4225 10535 4305
rect 10605 4225 10625 4305
rect 10695 4225 10715 4305
rect 10785 4225 10805 4305
rect 10875 4225 10895 4305
rect 10965 4225 10985 4305
rect 11055 4225 11075 4305
rect 11145 4225 11165 4305
rect 11235 4225 11255 4305
rect 11325 4225 11345 4305
rect 11415 4225 11435 4305
rect 11505 4225 11525 4305
rect 11595 4225 11615 4305
rect 11685 4225 11705 4305
rect 11775 4225 11795 4305
rect 11865 4225 11885 4305
rect 11955 4225 11975 4305
rect 12045 4225 12065 4305
rect 12135 4225 12155 4305
rect 12225 4225 12245 4305
rect 12315 4225 12335 4305
rect 12405 4225 12425 4305
rect 12495 4225 12515 4305
rect 12585 4225 12605 4305
rect 12675 4225 12695 4305
rect 12765 4225 12785 4305
rect 12855 4225 12875 4305
rect 12945 4225 12965 4305
rect 13035 4225 13055 4305
rect 13125 4225 13145 4305
rect 13215 4225 13235 4305
rect 13305 4225 13325 4305
rect 13395 4225 13415 4305
rect 13485 4225 13505 4305
rect 13575 4225 13595 4305
rect 13665 4225 13685 4305
rect 13755 4225 13775 4305
rect 13845 4225 13865 4305
rect 13935 4225 13955 4305
rect 14025 4225 14045 4305
rect 14115 4225 14135 4305
rect 14205 4225 14225 4305
rect 14295 4225 14315 4305
rect 14385 4225 14405 4305
rect 14475 4225 14495 4305
rect 14565 4225 14585 4305
rect 14655 4225 14675 4305
rect 14745 4225 14765 4305
rect 14835 4225 14855 4305
rect 14925 4225 14945 4305
rect 15015 4225 15035 4305
rect 15105 4225 15125 4305
rect 15195 4225 15215 4305
rect 15285 4225 15305 4305
rect 15375 4225 15395 4305
rect 15465 4225 15485 4305
rect 15555 4225 15575 4305
rect 15645 4225 15665 4305
rect 15735 4225 15755 4305
rect 15825 4225 15845 4305
rect 15915 4225 15935 4305
rect 16005 4225 16025 4305
rect 16095 4225 16115 4305
rect 16185 4225 16205 4305
rect 16275 4225 16295 4305
rect 16365 4225 16385 4305
rect 16455 4225 16475 4305
rect 16545 4225 16565 4305
rect 16635 4225 16655 4305
rect 16725 4225 16745 4305
rect 16815 4225 16835 4305
rect 16905 4225 16925 4305
rect 16995 4225 17015 4305
rect 17085 4225 17105 4305
rect 17175 4225 17195 4305
rect 17265 4225 17285 4305
rect 17355 4225 17375 4305
rect 17445 4225 17465 4305
rect 17535 4225 17555 4305
rect 17625 4225 17645 4305
rect 17715 4225 17735 4305
rect 17805 4225 17825 4305
rect 17895 4225 17915 4305
rect 17985 4225 18005 4305
rect 18075 4225 18095 4305
rect 18165 4225 18185 4305
rect 18255 4225 18275 4305
rect 18345 4225 18365 4305
rect 18435 4225 18455 4305
rect 18525 4225 18545 4305
rect 18615 4225 18635 4305
rect 18705 4225 18725 4305
rect 18795 4225 18815 4305
rect 18885 4225 18905 4305
rect 18975 4225 18995 4305
rect 19065 4225 19085 4305
rect 19155 4225 19175 4305
rect 19245 4225 19265 4305
rect 19335 4225 19355 4305
rect 19425 4225 19445 4305
rect 19515 4225 19535 4305
rect 19605 4225 19625 4305
rect 19695 4225 19715 4305
rect 19785 4225 19805 4305
rect 19875 4225 19895 4305
rect 19965 4225 19985 4305
rect 20685 4225 20705 4305
rect 10020 4170 10040 4190
rect 10200 4170 10220 4190
rect 10380 4170 10400 4190
rect 10560 4170 10580 4190
rect 10740 4170 10760 4190
rect 10920 4170 10940 4190
rect 11100 4170 11120 4190
rect 11280 4170 11300 4190
rect 11460 4170 11480 4190
rect 11640 4170 11660 4190
rect 11820 4170 11840 4190
rect 12000 4170 12020 4190
rect 12180 4170 12200 4190
rect 12360 4170 12380 4190
rect 12540 4170 12560 4190
rect 12720 4170 12740 4190
rect 12900 4170 12920 4190
rect 13080 4170 13100 4190
rect 13260 4170 13280 4190
rect 13440 4170 13460 4190
rect 13620 4170 13640 4190
rect 13800 4170 13820 4190
rect 13980 4170 14000 4190
rect 14160 4170 14180 4190
rect 14340 4170 14360 4190
rect 14520 4170 14540 4190
rect 14700 4170 14720 4190
rect 14880 4170 14900 4190
rect 15060 4170 15080 4190
rect 15240 4170 15260 4190
rect 15420 4170 15440 4190
rect 15600 4170 15620 4190
rect 15780 4170 15800 4190
rect 15960 4170 15980 4190
rect 16140 4170 16160 4190
rect 16320 4170 16340 4190
rect 16500 4170 16520 4190
rect 16680 4170 16700 4190
rect 16860 4170 16880 4190
rect 17040 4170 17060 4190
rect 17220 4170 17240 4190
rect 17400 4170 17420 4190
rect 17580 4170 17600 4190
rect 17760 4170 17780 4190
rect 17940 4170 17960 4190
rect 18120 4170 18140 4190
rect 18300 4170 18320 4190
rect 18480 4170 18500 4190
rect 18660 4170 18680 4190
rect 18840 4170 18860 4190
rect 19020 4170 19040 4190
rect 19200 4170 19220 4190
rect 19380 4170 19400 4190
rect 19560 4170 19580 4190
rect 19740 4170 19760 4190
rect 19920 4170 19940 4190
rect 9795 4085 9815 4105
rect 11370 4085 11390 4105
rect 11685 4085 11705 4105
rect 11910 4085 11930 4105
rect 12090 4085 12110 4105
rect 12630 4085 12650 4105
rect 20145 4085 20165 4105
rect 11460 4005 11480 4025
rect 12000 4005 12020 4025
rect 11640 3965 11660 3985
rect 11820 3965 11840 3985
rect 20325 3965 20345 3985
rect 10785 3925 10805 3945
rect 11145 3925 11165 3945
rect 12225 3925 12245 3945
rect 12585 3925 12605 3945
rect 20415 3925 20435 3945
rect 12270 3885 12290 3905
rect 12360 3885 12380 3905
rect 12405 3885 12425 3905
rect 12450 3885 12470 3905
rect 12540 3885 12560 3905
rect 20235 3885 20255 3905
rect 10920 3845 10940 3865
rect 11100 3845 11120 3865
rect 11550 3845 11570 3865
rect 11730 3845 11750 3865
rect 11505 3805 11525 3825
rect 11865 3805 11885 3825
rect 12045 3805 12065 3825
rect 10740 3765 10760 3785
rect 10965 3765 10985 3785
rect 11280 3765 11300 3785
rect 12180 3765 12200 3785
rect 12720 3765 12740 3785
rect 10830 3725 10850 3745
rect 11010 3725 11030 3745
rect 20505 3725 20525 3745
rect 10650 3685 10670 3705
rect 11190 3685 11210 3705
rect 20595 3685 20615 3705
rect 9930 3600 9950 3620
rect 10110 3600 10130 3620
rect 10290 3600 10310 3620
rect 10470 3600 10490 3620
rect 10650 3600 10670 3620
rect 10830 3600 10850 3620
rect 11010 3600 11030 3620
rect 11190 3600 11210 3620
rect 11370 3600 11390 3620
rect 11550 3600 11570 3620
rect 11730 3600 11750 3620
rect 11910 3600 11930 3620
rect 12090 3600 12110 3620
rect 12270 3600 12290 3620
rect 12450 3600 12470 3620
rect 12630 3600 12650 3620
rect 12810 3600 12830 3620
rect 12990 3600 13010 3620
rect 13170 3600 13190 3620
rect 13350 3600 13370 3620
rect 13530 3600 13550 3620
rect 13710 3600 13730 3620
rect 13890 3600 13910 3620
rect 14070 3600 14090 3620
rect 14250 3600 14270 3620
rect 14430 3600 14450 3620
rect 14610 3600 14630 3620
rect 14790 3600 14810 3620
rect 14970 3600 14990 3620
rect 15150 3600 15170 3620
rect 15330 3600 15350 3620
rect 15510 3600 15530 3620
rect 15690 3600 15710 3620
rect 15870 3600 15890 3620
rect 16050 3600 16070 3620
rect 16230 3600 16250 3620
rect 16410 3600 16430 3620
rect 16590 3600 16610 3620
rect 16770 3600 16790 3620
rect 16950 3600 16970 3620
rect 17130 3600 17150 3620
rect 17310 3600 17330 3620
rect 17490 3600 17510 3620
rect 17670 3600 17690 3620
rect 17850 3600 17870 3620
rect 18030 3600 18050 3620
rect 18210 3600 18230 3620
rect 18390 3600 18410 3620
rect 18570 3600 18590 3620
rect 18750 3600 18770 3620
rect 18930 3600 18950 3620
rect 19110 3600 19130 3620
rect 19290 3600 19310 3620
rect 19470 3600 19490 3620
rect 19650 3600 19670 3620
rect 19830 3600 19850 3620
rect 9165 3485 9185 3565
rect 9885 3485 9905 3565
rect 9975 3485 9995 3565
rect 10065 3485 10085 3565
rect 10155 3485 10175 3565
rect 10245 3485 10265 3565
rect 10335 3485 10355 3565
rect 10425 3485 10445 3565
rect 10515 3485 10535 3565
rect 10605 3485 10625 3565
rect 10695 3485 10715 3565
rect 10785 3485 10805 3565
rect 10875 3485 10895 3565
rect 10965 3485 10985 3565
rect 11055 3485 11075 3565
rect 11145 3485 11165 3565
rect 11235 3485 11255 3565
rect 11325 3485 11345 3565
rect 11415 3485 11435 3565
rect 11505 3485 11525 3565
rect 11595 3485 11615 3565
rect 11685 3485 11705 3565
rect 11775 3485 11795 3565
rect 11865 3485 11885 3565
rect 11955 3485 11975 3565
rect 12045 3485 12065 3565
rect 12135 3485 12155 3565
rect 12225 3485 12245 3565
rect 12315 3485 12335 3565
rect 12405 3485 12425 3565
rect 12495 3485 12515 3565
rect 12585 3485 12605 3565
rect 12675 3485 12695 3565
rect 12765 3485 12785 3565
rect 12855 3485 12875 3565
rect 12945 3485 12965 3565
rect 13035 3485 13055 3565
rect 13125 3485 13145 3565
rect 13215 3485 13235 3565
rect 13305 3485 13325 3565
rect 13395 3485 13415 3565
rect 13485 3485 13505 3565
rect 13575 3485 13595 3565
rect 13665 3485 13685 3565
rect 13755 3485 13775 3565
rect 13845 3485 13865 3565
rect 13935 3485 13955 3565
rect 14025 3485 14045 3565
rect 14115 3485 14135 3565
rect 14205 3485 14225 3565
rect 14295 3485 14315 3565
rect 14385 3485 14405 3565
rect 14475 3485 14495 3565
rect 14565 3485 14585 3565
rect 14655 3485 14675 3565
rect 14745 3485 14765 3565
rect 14835 3485 14855 3565
rect 14925 3485 14945 3565
rect 15015 3485 15035 3565
rect 15105 3485 15125 3565
rect 15195 3485 15215 3565
rect 15285 3485 15305 3565
rect 15375 3485 15395 3565
rect 15465 3485 15485 3565
rect 15555 3485 15575 3565
rect 15645 3485 15665 3565
rect 15735 3485 15755 3565
rect 15825 3485 15845 3565
rect 15915 3485 15935 3565
rect 16005 3485 16025 3565
rect 16095 3485 16115 3565
rect 16185 3485 16205 3565
rect 16275 3485 16295 3565
rect 16365 3485 16385 3565
rect 16455 3485 16475 3565
rect 16545 3485 16565 3565
rect 16635 3485 16655 3565
rect 16725 3485 16745 3565
rect 16815 3485 16835 3565
rect 16905 3485 16925 3565
rect 16995 3485 17015 3565
rect 17085 3485 17105 3565
rect 17175 3485 17195 3565
rect 17265 3485 17285 3565
rect 17355 3485 17375 3565
rect 17445 3485 17465 3565
rect 17535 3485 17555 3565
rect 17625 3485 17645 3565
rect 17715 3485 17735 3565
rect 17805 3485 17825 3565
rect 17895 3485 17915 3565
rect 17985 3485 18005 3565
rect 18075 3485 18095 3565
rect 18165 3485 18185 3565
rect 18255 3485 18275 3565
rect 18345 3485 18365 3565
rect 18435 3485 18455 3565
rect 18525 3485 18545 3565
rect 18615 3485 18635 3565
rect 18705 3485 18725 3565
rect 18795 3485 18815 3565
rect 18885 3485 18905 3565
rect 18975 3485 18995 3565
rect 19065 3485 19085 3565
rect 19155 3485 19175 3565
rect 19245 3485 19265 3565
rect 19335 3485 19355 3565
rect 19425 3485 19445 3565
rect 19515 3485 19535 3565
rect 19605 3485 19625 3565
rect 19695 3485 19715 3565
rect 19785 3485 19805 3565
rect 19875 3485 19895 3565
rect 19965 3485 19985 3565
rect 20685 3485 20705 3565
rect 9030 3425 9050 3445
rect 9165 3425 9185 3445
rect 9885 3425 9905 3445
rect 10065 3425 10085 3445
rect 10245 3425 10265 3445
rect 10425 3425 10445 3445
rect 10605 3425 10625 3445
rect 10785 3425 10805 3445
rect 10965 3425 10985 3445
rect 11145 3425 11165 3445
rect 11325 3425 11345 3445
rect 11505 3425 11525 3445
rect 11685 3425 11705 3445
rect 11865 3425 11885 3445
rect 12045 3425 12065 3445
rect 12225 3425 12245 3445
rect 12405 3425 12425 3445
rect 12585 3425 12605 3445
rect 12765 3425 12785 3445
rect 12945 3425 12965 3445
rect 13125 3425 13145 3445
rect 13305 3425 13325 3445
rect 13485 3425 13505 3445
rect 13665 3425 13685 3445
rect 13845 3425 13865 3445
rect 14025 3425 14045 3445
rect 14205 3425 14225 3445
rect 14385 3425 14405 3445
rect 14565 3425 14585 3445
rect 14745 3425 14765 3445
rect 14925 3425 14945 3445
rect 15105 3425 15125 3445
rect 15285 3425 15305 3445
rect 15465 3425 15485 3445
rect 15645 3425 15665 3445
rect 15825 3425 15845 3445
rect 16005 3425 16025 3445
rect 16185 3425 16205 3445
rect 16365 3425 16385 3445
rect 16545 3425 16565 3445
rect 16725 3425 16745 3445
rect 16905 3425 16925 3445
rect 17085 3425 17105 3445
rect 17265 3425 17285 3445
rect 17445 3425 17465 3445
rect 17625 3425 17645 3445
rect 17805 3425 17825 3445
rect 17985 3425 18005 3445
rect 18165 3425 18185 3445
rect 18345 3425 18365 3445
rect 18525 3425 18545 3445
rect 18705 3425 18725 3445
rect 18885 3425 18905 3445
rect 19065 3425 19085 3445
rect 19245 3425 19265 3445
rect 19425 3425 19445 3445
rect 19605 3425 19625 3445
rect 19785 3425 19805 3445
rect 19965 3425 19985 3445
rect 20685 3425 20705 3445
rect 20820 3425 20840 3445
<< metal1 >>
rect 9020 3450 9060 4375
rect 9155 4370 9195 4375
rect 9155 4340 9160 4370
rect 9190 4340 9195 4370
rect 9155 4335 9195 4340
rect 9165 4315 9185 4335
rect 9255 4315 9275 4375
rect 9345 4315 9365 4375
rect 9435 4315 9455 4375
rect 9525 4315 9545 4375
rect 9615 4315 9635 4375
rect 9705 4315 9725 4375
rect 9795 4315 9815 4375
rect 9875 4370 9915 4375
rect 9875 4340 9880 4370
rect 9910 4340 9915 4370
rect 9875 4335 9915 4340
rect 10055 4370 10095 4375
rect 10055 4340 10060 4370
rect 10090 4340 10095 4370
rect 10055 4335 10095 4340
rect 10235 4370 10275 4375
rect 10235 4340 10240 4370
rect 10270 4340 10275 4370
rect 10235 4335 10275 4340
rect 10415 4370 10455 4375
rect 10415 4340 10420 4370
rect 10450 4340 10455 4370
rect 10415 4335 10455 4340
rect 10595 4370 10635 4375
rect 10595 4340 10600 4370
rect 10630 4340 10635 4370
rect 10595 4335 10635 4340
rect 10775 4370 10815 4375
rect 10775 4340 10780 4370
rect 10810 4340 10815 4370
rect 10775 4335 10815 4340
rect 10955 4370 10995 4375
rect 10955 4340 10960 4370
rect 10990 4340 10995 4370
rect 10955 4335 10995 4340
rect 11135 4370 11175 4375
rect 11135 4340 11140 4370
rect 11170 4340 11175 4370
rect 11135 4335 11175 4340
rect 11315 4370 11355 4375
rect 11315 4340 11320 4370
rect 11350 4340 11355 4370
rect 11315 4335 11355 4340
rect 11495 4370 11535 4375
rect 11495 4340 11500 4370
rect 11530 4340 11535 4370
rect 11495 4335 11535 4340
rect 11675 4370 11715 4375
rect 11675 4340 11680 4370
rect 11710 4340 11715 4370
rect 11675 4335 11715 4340
rect 11855 4370 11895 4375
rect 11855 4340 11860 4370
rect 11890 4340 11895 4370
rect 11855 4335 11895 4340
rect 12035 4370 12075 4375
rect 12035 4340 12040 4370
rect 12070 4340 12075 4370
rect 12035 4335 12075 4340
rect 12215 4370 12255 4375
rect 12215 4340 12220 4370
rect 12250 4340 12255 4370
rect 12215 4335 12255 4340
rect 12395 4370 12435 4375
rect 12395 4340 12400 4370
rect 12430 4340 12435 4370
rect 12395 4335 12435 4340
rect 12575 4370 12615 4375
rect 12575 4340 12580 4370
rect 12610 4340 12615 4370
rect 12575 4335 12615 4340
rect 12755 4370 12795 4375
rect 12755 4340 12760 4370
rect 12790 4340 12795 4370
rect 12755 4335 12795 4340
rect 12935 4370 12975 4375
rect 12935 4340 12940 4370
rect 12970 4340 12975 4370
rect 12935 4335 12975 4340
rect 13115 4370 13155 4375
rect 13115 4340 13120 4370
rect 13150 4340 13155 4370
rect 13115 4335 13155 4340
rect 13295 4370 13335 4375
rect 13295 4340 13300 4370
rect 13330 4340 13335 4370
rect 13295 4335 13335 4340
rect 13475 4370 13515 4375
rect 13475 4340 13480 4370
rect 13510 4340 13515 4370
rect 13475 4335 13515 4340
rect 13655 4370 13695 4375
rect 13655 4340 13660 4370
rect 13690 4340 13695 4370
rect 13655 4335 13695 4340
rect 13835 4370 13875 4375
rect 13835 4340 13840 4370
rect 13870 4340 13875 4370
rect 13835 4335 13875 4340
rect 14015 4370 14055 4375
rect 14015 4340 14020 4370
rect 14050 4340 14055 4370
rect 14015 4335 14055 4340
rect 14195 4370 14235 4375
rect 14195 4340 14200 4370
rect 14230 4340 14235 4370
rect 14195 4335 14235 4340
rect 14375 4370 14415 4375
rect 14375 4340 14380 4370
rect 14410 4340 14415 4370
rect 14375 4335 14415 4340
rect 14555 4370 14595 4375
rect 14555 4340 14560 4370
rect 14590 4340 14595 4370
rect 14555 4335 14595 4340
rect 14735 4370 14775 4375
rect 14735 4340 14740 4370
rect 14770 4340 14775 4370
rect 14735 4335 14775 4340
rect 14915 4370 14955 4375
rect 14915 4340 14920 4370
rect 14950 4340 14955 4370
rect 14915 4335 14955 4340
rect 15095 4370 15135 4375
rect 15095 4340 15100 4370
rect 15130 4340 15135 4370
rect 15095 4335 15135 4340
rect 15275 4370 15315 4375
rect 15275 4340 15280 4370
rect 15310 4340 15315 4370
rect 15275 4335 15315 4340
rect 15455 4370 15495 4375
rect 15455 4340 15460 4370
rect 15490 4340 15495 4370
rect 15455 4335 15495 4340
rect 15635 4370 15675 4375
rect 15635 4340 15640 4370
rect 15670 4340 15675 4370
rect 15635 4335 15675 4340
rect 15815 4370 15855 4375
rect 15815 4340 15820 4370
rect 15850 4340 15855 4370
rect 15815 4335 15855 4340
rect 15995 4370 16035 4375
rect 15995 4340 16000 4370
rect 16030 4340 16035 4370
rect 15995 4335 16035 4340
rect 16175 4370 16215 4375
rect 16175 4340 16180 4370
rect 16210 4340 16215 4370
rect 16175 4335 16215 4340
rect 16355 4370 16395 4375
rect 16355 4340 16360 4370
rect 16390 4340 16395 4370
rect 16355 4335 16395 4340
rect 16535 4370 16575 4375
rect 16535 4340 16540 4370
rect 16570 4340 16575 4370
rect 16535 4335 16575 4340
rect 16715 4370 16755 4375
rect 16715 4340 16720 4370
rect 16750 4340 16755 4370
rect 16715 4335 16755 4340
rect 16895 4370 16935 4375
rect 16895 4340 16900 4370
rect 16930 4340 16935 4370
rect 16895 4335 16935 4340
rect 17075 4370 17115 4375
rect 17075 4340 17080 4370
rect 17110 4340 17115 4370
rect 17075 4335 17115 4340
rect 17255 4370 17295 4375
rect 17255 4340 17260 4370
rect 17290 4340 17295 4370
rect 17255 4335 17295 4340
rect 17435 4370 17475 4375
rect 17435 4340 17440 4370
rect 17470 4340 17475 4370
rect 17435 4335 17475 4340
rect 17615 4370 17655 4375
rect 17615 4340 17620 4370
rect 17650 4340 17655 4370
rect 17615 4335 17655 4340
rect 17795 4370 17835 4375
rect 17795 4340 17800 4370
rect 17830 4340 17835 4370
rect 17795 4335 17835 4340
rect 17975 4370 18015 4375
rect 17975 4340 17980 4370
rect 18010 4340 18015 4370
rect 17975 4335 18015 4340
rect 18155 4370 18195 4375
rect 18155 4340 18160 4370
rect 18190 4340 18195 4370
rect 18155 4335 18195 4340
rect 18335 4370 18375 4375
rect 18335 4340 18340 4370
rect 18370 4340 18375 4370
rect 18335 4335 18375 4340
rect 18515 4370 18555 4375
rect 18515 4340 18520 4370
rect 18550 4340 18555 4370
rect 18515 4335 18555 4340
rect 18695 4370 18735 4375
rect 18695 4340 18700 4370
rect 18730 4340 18735 4370
rect 18695 4335 18735 4340
rect 18875 4370 18915 4375
rect 18875 4340 18880 4370
rect 18910 4340 18915 4370
rect 18875 4335 18915 4340
rect 19055 4370 19095 4375
rect 19055 4340 19060 4370
rect 19090 4340 19095 4370
rect 19055 4335 19095 4340
rect 19235 4370 19275 4375
rect 19235 4340 19240 4370
rect 19270 4340 19275 4370
rect 19235 4335 19275 4340
rect 19415 4370 19455 4375
rect 19415 4340 19420 4370
rect 19450 4340 19455 4370
rect 19415 4335 19455 4340
rect 19595 4370 19635 4375
rect 19595 4340 19600 4370
rect 19630 4340 19635 4370
rect 19595 4335 19635 4340
rect 19775 4370 19815 4375
rect 19775 4340 19780 4370
rect 19810 4340 19815 4370
rect 19775 4335 19815 4340
rect 19955 4370 19995 4375
rect 19955 4340 19960 4370
rect 19990 4340 19995 4370
rect 19955 4335 19995 4340
rect 9885 4315 9905 4335
rect 10605 4315 10625 4335
rect 11325 4315 11345 4335
rect 12045 4315 12065 4335
rect 12765 4315 12785 4335
rect 14925 4315 14945 4335
rect 17085 4315 17105 4335
rect 19245 4315 19265 4335
rect 19425 4315 19445 4335
rect 19605 4315 19625 4335
rect 19785 4315 19805 4335
rect 19965 4315 19985 4335
rect 20055 4315 20075 4375
rect 20145 4315 20165 4375
rect 20235 4315 20255 4375
rect 20325 4315 20345 4375
rect 20415 4315 20435 4375
rect 20505 4315 20525 4375
rect 20595 4315 20615 4375
rect 20675 4370 20715 4375
rect 20675 4340 20680 4370
rect 20710 4340 20715 4370
rect 20675 4335 20715 4340
rect 20685 4315 20705 4335
rect 9160 4305 9190 4315
rect 9160 4225 9165 4305
rect 9185 4225 9190 4305
rect 9160 4215 9190 4225
rect 9250 4215 9280 4315
rect 9340 4215 9370 4315
rect 9430 4215 9460 4315
rect 9520 4215 9550 4315
rect 9610 4215 9640 4315
rect 9700 4215 9730 4315
rect 9790 4215 9820 4315
rect 9880 4305 9910 4315
rect 9880 4225 9885 4305
rect 9905 4225 9910 4305
rect 9880 4215 9910 4225
rect 9970 4305 10000 4315
rect 9970 4225 9975 4305
rect 9995 4225 10000 4305
rect 9970 4215 10000 4225
rect 10060 4305 10090 4315
rect 10060 4225 10065 4305
rect 10085 4225 10090 4305
rect 10060 4215 10090 4225
rect 10150 4305 10180 4315
rect 10150 4225 10155 4305
rect 10175 4225 10180 4305
rect 10150 4215 10180 4225
rect 10240 4305 10270 4315
rect 10240 4225 10245 4305
rect 10265 4225 10270 4305
rect 10240 4215 10270 4225
rect 10330 4305 10360 4315
rect 10330 4225 10335 4305
rect 10355 4225 10360 4305
rect 10330 4215 10360 4225
rect 10420 4305 10450 4315
rect 10420 4225 10425 4305
rect 10445 4225 10450 4305
rect 10420 4215 10450 4225
rect 10510 4305 10540 4315
rect 10510 4225 10515 4305
rect 10535 4225 10540 4305
rect 10510 4215 10540 4225
rect 10600 4305 10630 4315
rect 10600 4225 10605 4305
rect 10625 4225 10630 4305
rect 10600 4215 10630 4225
rect 10690 4305 10720 4315
rect 10690 4225 10695 4305
rect 10715 4225 10720 4305
rect 10690 4215 10720 4225
rect 10780 4305 10810 4315
rect 10780 4225 10785 4305
rect 10805 4225 10810 4305
rect 10780 4215 10810 4225
rect 10870 4305 10900 4315
rect 10870 4225 10875 4305
rect 10895 4225 10900 4305
rect 10870 4215 10900 4225
rect 10960 4305 10990 4315
rect 10960 4225 10965 4305
rect 10985 4225 10990 4305
rect 10960 4215 10990 4225
rect 11050 4305 11080 4315
rect 11050 4225 11055 4305
rect 11075 4225 11080 4305
rect 11050 4215 11080 4225
rect 11140 4305 11170 4315
rect 11140 4225 11145 4305
rect 11165 4225 11170 4305
rect 11140 4215 11170 4225
rect 11230 4305 11260 4315
rect 11230 4225 11235 4305
rect 11255 4225 11260 4305
rect 11230 4215 11260 4225
rect 11320 4305 11350 4315
rect 11320 4225 11325 4305
rect 11345 4225 11350 4305
rect 11320 4215 11350 4225
rect 11410 4305 11440 4315
rect 11410 4225 11415 4305
rect 11435 4225 11440 4305
rect 11410 4215 11440 4225
rect 11500 4305 11530 4315
rect 11500 4225 11505 4305
rect 11525 4225 11530 4305
rect 11500 4215 11530 4225
rect 11590 4305 11620 4315
rect 11590 4225 11595 4305
rect 11615 4225 11620 4305
rect 11590 4215 11620 4225
rect 11680 4305 11710 4315
rect 11680 4225 11685 4305
rect 11705 4225 11710 4305
rect 11680 4215 11710 4225
rect 11770 4305 11800 4315
rect 11770 4225 11775 4305
rect 11795 4225 11800 4305
rect 11770 4215 11800 4225
rect 11860 4305 11890 4315
rect 11860 4225 11865 4305
rect 11885 4225 11890 4305
rect 11860 4215 11890 4225
rect 11950 4305 11980 4315
rect 11950 4225 11955 4305
rect 11975 4225 11980 4305
rect 11950 4215 11980 4225
rect 12040 4305 12070 4315
rect 12040 4225 12045 4305
rect 12065 4225 12070 4305
rect 12040 4215 12070 4225
rect 12130 4305 12160 4315
rect 12130 4225 12135 4305
rect 12155 4225 12160 4305
rect 12130 4215 12160 4225
rect 12220 4305 12250 4315
rect 12220 4225 12225 4305
rect 12245 4225 12250 4305
rect 12220 4215 12250 4225
rect 12310 4305 12340 4315
rect 12310 4225 12315 4305
rect 12335 4225 12340 4305
rect 12310 4215 12340 4225
rect 12400 4305 12430 4315
rect 12400 4225 12405 4305
rect 12425 4225 12430 4305
rect 12400 4215 12430 4225
rect 12490 4305 12520 4315
rect 12490 4225 12495 4305
rect 12515 4225 12520 4305
rect 12490 4215 12520 4225
rect 12580 4305 12610 4315
rect 12580 4225 12585 4305
rect 12605 4225 12610 4305
rect 12580 4215 12610 4225
rect 12670 4305 12700 4315
rect 12670 4225 12675 4305
rect 12695 4225 12700 4305
rect 12670 4215 12700 4225
rect 12760 4305 12790 4315
rect 12760 4225 12765 4305
rect 12785 4225 12790 4305
rect 12760 4215 12790 4225
rect 12850 4305 12880 4315
rect 12850 4225 12855 4305
rect 12875 4225 12880 4305
rect 12850 4215 12880 4225
rect 12940 4305 12970 4315
rect 12940 4225 12945 4305
rect 12965 4225 12970 4305
rect 12940 4215 12970 4225
rect 13030 4305 13060 4315
rect 13030 4225 13035 4305
rect 13055 4225 13060 4305
rect 13030 4215 13060 4225
rect 13120 4305 13150 4315
rect 13120 4225 13125 4305
rect 13145 4225 13150 4305
rect 13120 4215 13150 4225
rect 13210 4305 13240 4315
rect 13210 4225 13215 4305
rect 13235 4225 13240 4305
rect 13210 4215 13240 4225
rect 13300 4305 13330 4315
rect 13300 4225 13305 4305
rect 13325 4225 13330 4305
rect 13300 4215 13330 4225
rect 13390 4305 13420 4315
rect 13390 4225 13395 4305
rect 13415 4225 13420 4305
rect 13390 4215 13420 4225
rect 13480 4305 13510 4315
rect 13480 4225 13485 4305
rect 13505 4225 13510 4305
rect 13480 4215 13510 4225
rect 13570 4305 13600 4315
rect 13570 4225 13575 4305
rect 13595 4225 13600 4305
rect 13570 4215 13600 4225
rect 13660 4305 13690 4315
rect 13660 4225 13665 4305
rect 13685 4225 13690 4305
rect 13660 4215 13690 4225
rect 13750 4305 13780 4315
rect 13750 4225 13755 4305
rect 13775 4225 13780 4305
rect 13750 4215 13780 4225
rect 13840 4305 13870 4315
rect 13840 4225 13845 4305
rect 13865 4225 13870 4305
rect 13840 4215 13870 4225
rect 13930 4305 13960 4315
rect 13930 4225 13935 4305
rect 13955 4225 13960 4305
rect 13930 4215 13960 4225
rect 14020 4305 14050 4315
rect 14020 4225 14025 4305
rect 14045 4225 14050 4305
rect 14020 4215 14050 4225
rect 14110 4305 14140 4315
rect 14110 4225 14115 4305
rect 14135 4225 14140 4305
rect 14110 4215 14140 4225
rect 14200 4305 14230 4315
rect 14200 4225 14205 4305
rect 14225 4225 14230 4305
rect 14200 4215 14230 4225
rect 14290 4305 14320 4315
rect 14290 4225 14295 4305
rect 14315 4225 14320 4305
rect 14290 4215 14320 4225
rect 14380 4305 14410 4315
rect 14380 4225 14385 4305
rect 14405 4225 14410 4305
rect 14380 4215 14410 4225
rect 14470 4305 14500 4315
rect 14470 4225 14475 4305
rect 14495 4225 14500 4305
rect 14470 4215 14500 4225
rect 14560 4305 14590 4315
rect 14560 4225 14565 4305
rect 14585 4225 14590 4305
rect 14560 4215 14590 4225
rect 14650 4305 14680 4315
rect 14650 4225 14655 4305
rect 14675 4225 14680 4305
rect 14650 4215 14680 4225
rect 14740 4305 14770 4315
rect 14740 4225 14745 4305
rect 14765 4225 14770 4305
rect 14740 4215 14770 4225
rect 14830 4305 14860 4315
rect 14830 4225 14835 4305
rect 14855 4225 14860 4305
rect 14830 4215 14860 4225
rect 14920 4305 14950 4315
rect 14920 4225 14925 4305
rect 14945 4225 14950 4305
rect 14920 4215 14950 4225
rect 15010 4305 15040 4315
rect 15010 4225 15015 4305
rect 15035 4225 15040 4305
rect 15010 4215 15040 4225
rect 15100 4305 15130 4315
rect 15100 4225 15105 4305
rect 15125 4225 15130 4305
rect 15100 4215 15130 4225
rect 15190 4305 15220 4315
rect 15190 4225 15195 4305
rect 15215 4225 15220 4305
rect 15190 4215 15220 4225
rect 15280 4305 15310 4315
rect 15280 4225 15285 4305
rect 15305 4225 15310 4305
rect 15280 4215 15310 4225
rect 15370 4305 15400 4315
rect 15370 4225 15375 4305
rect 15395 4225 15400 4305
rect 15370 4215 15400 4225
rect 15460 4305 15490 4315
rect 15460 4225 15465 4305
rect 15485 4225 15490 4305
rect 15460 4215 15490 4225
rect 15550 4305 15580 4315
rect 15550 4225 15555 4305
rect 15575 4225 15580 4305
rect 15550 4215 15580 4225
rect 15640 4305 15670 4315
rect 15640 4225 15645 4305
rect 15665 4225 15670 4305
rect 15640 4215 15670 4225
rect 15730 4305 15760 4315
rect 15730 4225 15735 4305
rect 15755 4225 15760 4305
rect 15730 4215 15760 4225
rect 15820 4305 15850 4315
rect 15820 4225 15825 4305
rect 15845 4225 15850 4305
rect 15820 4215 15850 4225
rect 15910 4305 15940 4315
rect 15910 4225 15915 4305
rect 15935 4225 15940 4305
rect 15910 4215 15940 4225
rect 16000 4305 16030 4315
rect 16000 4225 16005 4305
rect 16025 4225 16030 4305
rect 16000 4215 16030 4225
rect 16090 4305 16120 4315
rect 16090 4225 16095 4305
rect 16115 4225 16120 4305
rect 16090 4215 16120 4225
rect 16180 4305 16210 4315
rect 16180 4225 16185 4305
rect 16205 4225 16210 4305
rect 16180 4215 16210 4225
rect 16270 4305 16300 4315
rect 16270 4225 16275 4305
rect 16295 4225 16300 4305
rect 16270 4215 16300 4225
rect 16360 4305 16390 4315
rect 16360 4225 16365 4305
rect 16385 4225 16390 4305
rect 16360 4215 16390 4225
rect 16450 4305 16480 4315
rect 16450 4225 16455 4305
rect 16475 4225 16480 4305
rect 16450 4215 16480 4225
rect 16540 4305 16570 4315
rect 16540 4225 16545 4305
rect 16565 4225 16570 4305
rect 16540 4215 16570 4225
rect 16630 4305 16660 4315
rect 16630 4225 16635 4305
rect 16655 4225 16660 4305
rect 16630 4215 16660 4225
rect 16720 4305 16750 4315
rect 16720 4225 16725 4305
rect 16745 4225 16750 4305
rect 16720 4215 16750 4225
rect 16810 4305 16840 4315
rect 16810 4225 16815 4305
rect 16835 4225 16840 4305
rect 16810 4215 16840 4225
rect 16900 4305 16930 4315
rect 16900 4225 16905 4305
rect 16925 4225 16930 4305
rect 16900 4215 16930 4225
rect 16990 4305 17020 4315
rect 16990 4225 16995 4305
rect 17015 4225 17020 4305
rect 16990 4215 17020 4225
rect 17080 4305 17110 4315
rect 17080 4225 17085 4305
rect 17105 4225 17110 4305
rect 17080 4215 17110 4225
rect 17170 4305 17200 4315
rect 17170 4225 17175 4305
rect 17195 4225 17200 4305
rect 17170 4215 17200 4225
rect 17260 4305 17290 4315
rect 17260 4225 17265 4305
rect 17285 4225 17290 4305
rect 17260 4215 17290 4225
rect 17350 4305 17380 4315
rect 17350 4225 17355 4305
rect 17375 4225 17380 4305
rect 17350 4215 17380 4225
rect 17440 4305 17470 4315
rect 17440 4225 17445 4305
rect 17465 4225 17470 4305
rect 17440 4215 17470 4225
rect 17530 4305 17560 4315
rect 17530 4225 17535 4305
rect 17555 4225 17560 4305
rect 17530 4215 17560 4225
rect 17620 4305 17650 4315
rect 17620 4225 17625 4305
rect 17645 4225 17650 4305
rect 17620 4215 17650 4225
rect 17710 4305 17740 4315
rect 17710 4225 17715 4305
rect 17735 4225 17740 4305
rect 17710 4215 17740 4225
rect 17800 4305 17830 4315
rect 17800 4225 17805 4305
rect 17825 4225 17830 4305
rect 17800 4215 17830 4225
rect 17890 4305 17920 4315
rect 17890 4225 17895 4305
rect 17915 4225 17920 4305
rect 17890 4215 17920 4225
rect 17980 4305 18010 4315
rect 17980 4225 17985 4305
rect 18005 4225 18010 4305
rect 17980 4215 18010 4225
rect 18070 4305 18100 4315
rect 18070 4225 18075 4305
rect 18095 4225 18100 4305
rect 18070 4215 18100 4225
rect 18160 4305 18190 4315
rect 18160 4225 18165 4305
rect 18185 4225 18190 4305
rect 18160 4215 18190 4225
rect 18250 4305 18280 4315
rect 18250 4225 18255 4305
rect 18275 4225 18280 4305
rect 18250 4215 18280 4225
rect 18340 4305 18370 4315
rect 18340 4225 18345 4305
rect 18365 4225 18370 4305
rect 18340 4215 18370 4225
rect 18430 4305 18460 4315
rect 18430 4225 18435 4305
rect 18455 4225 18460 4305
rect 18430 4215 18460 4225
rect 18520 4305 18550 4315
rect 18520 4225 18525 4305
rect 18545 4225 18550 4305
rect 18520 4215 18550 4225
rect 18610 4305 18640 4315
rect 18610 4225 18615 4305
rect 18635 4225 18640 4305
rect 18610 4215 18640 4225
rect 18700 4305 18730 4315
rect 18700 4225 18705 4305
rect 18725 4225 18730 4305
rect 18700 4215 18730 4225
rect 18790 4305 18820 4315
rect 18790 4225 18795 4305
rect 18815 4225 18820 4305
rect 18790 4215 18820 4225
rect 18880 4305 18910 4315
rect 18880 4225 18885 4305
rect 18905 4225 18910 4305
rect 18880 4215 18910 4225
rect 18970 4305 19000 4315
rect 18970 4225 18975 4305
rect 18995 4225 19000 4305
rect 18970 4215 19000 4225
rect 19060 4305 19090 4315
rect 19060 4225 19065 4305
rect 19085 4225 19090 4305
rect 19060 4215 19090 4225
rect 19150 4305 19180 4315
rect 19150 4225 19155 4305
rect 19175 4225 19180 4305
rect 19150 4215 19180 4225
rect 19240 4305 19270 4315
rect 19240 4225 19245 4305
rect 19265 4225 19270 4305
rect 19240 4215 19270 4225
rect 19330 4305 19360 4315
rect 19330 4225 19335 4305
rect 19355 4225 19360 4305
rect 19330 4215 19360 4225
rect 19420 4305 19450 4315
rect 19420 4225 19425 4305
rect 19445 4225 19450 4305
rect 19420 4215 19450 4225
rect 19510 4305 19540 4315
rect 19510 4225 19515 4305
rect 19535 4225 19540 4305
rect 19510 4215 19540 4225
rect 19600 4305 19630 4315
rect 19600 4225 19605 4305
rect 19625 4225 19630 4305
rect 19600 4215 19630 4225
rect 19690 4305 19720 4315
rect 19690 4225 19695 4305
rect 19715 4225 19720 4305
rect 19690 4215 19720 4225
rect 19780 4305 19810 4315
rect 19780 4225 19785 4305
rect 19805 4225 19810 4305
rect 19780 4215 19810 4225
rect 19870 4305 19900 4315
rect 19870 4225 19875 4305
rect 19895 4225 19900 4305
rect 19870 4215 19900 4225
rect 19960 4305 19990 4315
rect 19960 4225 19965 4305
rect 19985 4225 19990 4305
rect 19960 4215 19990 4225
rect 20050 4215 20080 4315
rect 20140 4215 20170 4315
rect 20230 4215 20260 4315
rect 20320 4215 20350 4315
rect 20410 4215 20440 4315
rect 20500 4215 20530 4315
rect 20590 4215 20620 4315
rect 20680 4305 20710 4315
rect 20680 4225 20685 4305
rect 20705 4225 20710 4305
rect 20680 4215 20710 4225
rect 9255 3575 9275 4215
rect 9345 3575 9365 4215
rect 9435 3575 9455 4215
rect 9525 3575 9545 4215
rect 9615 3575 9635 4215
rect 9705 3575 9725 4215
rect 9795 4110 9815 4215
rect 10020 4195 10040 4200
rect 10200 4195 10220 4200
rect 10380 4195 10400 4200
rect 10560 4195 10580 4200
rect 10740 4195 10760 4200
rect 10015 4190 10045 4195
rect 10015 4170 10020 4190
rect 10040 4170 10045 4190
rect 10015 4165 10045 4170
rect 10195 4190 10225 4195
rect 10195 4170 10200 4190
rect 10220 4170 10225 4190
rect 10195 4165 10225 4170
rect 10375 4190 10405 4195
rect 10375 4170 10380 4190
rect 10400 4170 10405 4190
rect 10375 4165 10405 4170
rect 10555 4190 10585 4195
rect 10555 4170 10560 4190
rect 10580 4170 10585 4190
rect 10555 4165 10585 4170
rect 10735 4190 10765 4195
rect 10735 4170 10740 4190
rect 10760 4170 10765 4190
rect 10735 4165 10765 4170
rect 10020 4160 10040 4165
rect 10200 4160 10220 4165
rect 10380 4160 10400 4165
rect 10560 4160 10580 4165
rect 9790 4105 9820 4110
rect 9790 4085 9795 4105
rect 9815 4085 9820 4105
rect 9790 4080 9820 4085
rect 9795 3575 9815 4080
rect 10740 3790 10760 4165
rect 10785 3950 10805 4215
rect 10920 4195 10940 4200
rect 10915 4190 10945 4195
rect 10915 4170 10920 4190
rect 10940 4170 10945 4190
rect 10915 4165 10945 4170
rect 10780 3945 10810 3950
rect 10780 3925 10785 3945
rect 10805 3925 10810 3945
rect 10780 3920 10810 3925
rect 10785 3915 10805 3920
rect 10920 3870 10940 4165
rect 10915 3865 10945 3870
rect 10915 3845 10920 3865
rect 10940 3845 10945 3865
rect 10915 3840 10945 3845
rect 10920 3835 10940 3840
rect 10965 3790 10985 4215
rect 11100 4195 11120 4200
rect 11095 4190 11125 4195
rect 11095 4170 11100 4190
rect 11120 4170 11125 4190
rect 11095 4165 11125 4170
rect 11100 3870 11120 4165
rect 11145 3950 11165 4215
rect 11280 4195 11300 4200
rect 11460 4195 11480 4200
rect 11640 4195 11660 4200
rect 11275 4190 11305 4195
rect 11275 4170 11280 4190
rect 11300 4170 11305 4190
rect 11275 4165 11305 4170
rect 11455 4190 11485 4195
rect 11455 4170 11460 4190
rect 11480 4170 11485 4190
rect 11455 4165 11485 4170
rect 11635 4190 11665 4195
rect 11635 4170 11640 4190
rect 11660 4170 11665 4190
rect 11635 4165 11665 4170
rect 11140 3945 11170 3950
rect 11140 3925 11145 3945
rect 11165 3925 11170 3945
rect 11140 3920 11170 3925
rect 11145 3915 11165 3920
rect 11095 3865 11125 3870
rect 11095 3845 11100 3865
rect 11120 3845 11125 3865
rect 11095 3840 11125 3845
rect 11100 3835 11120 3840
rect 11280 3790 11300 4165
rect 11370 4110 11390 4115
rect 11365 4105 11395 4110
rect 11365 4085 11370 4105
rect 11390 4085 11395 4105
rect 11365 4080 11395 4085
rect 10735 3785 10765 3790
rect 10735 3765 10740 3785
rect 10760 3765 10765 3785
rect 10735 3760 10765 3765
rect 10960 3785 10990 3790
rect 10960 3765 10965 3785
rect 10985 3765 10990 3785
rect 10960 3760 10990 3765
rect 11275 3785 11305 3790
rect 11275 3765 11280 3785
rect 11300 3765 11305 3785
rect 11275 3760 11305 3765
rect 10740 3755 10760 3760
rect 10830 3750 10850 3755
rect 10825 3745 10855 3750
rect 10825 3725 10830 3745
rect 10850 3725 10855 3745
rect 10825 3720 10855 3725
rect 10650 3710 10670 3715
rect 10645 3705 10675 3710
rect 10645 3685 10650 3705
rect 10670 3685 10675 3705
rect 10645 3680 10675 3685
rect 9930 3625 9950 3630
rect 10110 3625 10130 3630
rect 10290 3625 10310 3630
rect 10470 3625 10490 3630
rect 10650 3625 10670 3680
rect 10830 3625 10850 3720
rect 9925 3620 9955 3625
rect 9925 3600 9930 3620
rect 9950 3600 9955 3620
rect 9925 3595 9955 3600
rect 10105 3620 10135 3625
rect 10105 3600 10110 3620
rect 10130 3600 10135 3620
rect 10105 3595 10135 3600
rect 10285 3620 10315 3625
rect 10285 3600 10290 3620
rect 10310 3600 10315 3620
rect 10285 3595 10315 3600
rect 10465 3620 10495 3625
rect 10465 3600 10470 3620
rect 10490 3600 10495 3620
rect 10465 3595 10495 3600
rect 10645 3620 10675 3625
rect 10645 3600 10650 3620
rect 10670 3600 10675 3620
rect 10645 3595 10675 3600
rect 10825 3620 10855 3625
rect 10825 3600 10830 3620
rect 10850 3600 10855 3620
rect 10825 3595 10855 3600
rect 9930 3590 9950 3595
rect 10110 3590 10130 3595
rect 10290 3590 10310 3595
rect 10470 3590 10490 3595
rect 10650 3590 10670 3595
rect 10830 3590 10850 3595
rect 10605 3575 10625 3580
rect 10965 3575 10985 3760
rect 11280 3755 11300 3760
rect 11010 3750 11030 3755
rect 11005 3745 11035 3750
rect 11005 3725 11010 3745
rect 11030 3725 11035 3745
rect 11005 3720 11035 3725
rect 11010 3625 11030 3720
rect 11190 3710 11210 3715
rect 11185 3705 11215 3710
rect 11185 3685 11190 3705
rect 11210 3685 11215 3705
rect 11185 3680 11215 3685
rect 11190 3625 11210 3680
rect 11370 3625 11390 4080
rect 11460 4030 11480 4165
rect 11455 4025 11485 4030
rect 11455 4005 11460 4025
rect 11480 4005 11485 4025
rect 11455 4000 11485 4005
rect 11460 3995 11480 4000
rect 11640 3990 11660 4165
rect 11685 4110 11705 4215
rect 11865 4210 11885 4215
rect 11820 4195 11840 4200
rect 12000 4195 12020 4200
rect 12180 4195 12200 4200
rect 11815 4190 11845 4195
rect 11815 4170 11820 4190
rect 11840 4170 11845 4190
rect 11815 4165 11845 4170
rect 11995 4190 12025 4195
rect 11995 4170 12000 4190
rect 12020 4170 12025 4190
rect 11995 4165 12025 4170
rect 12175 4190 12205 4195
rect 12175 4170 12180 4190
rect 12200 4170 12205 4190
rect 12175 4165 12205 4170
rect 11680 4105 11710 4110
rect 11680 4085 11685 4105
rect 11705 4085 11710 4105
rect 11680 4080 11710 4085
rect 11635 3985 11665 3990
rect 11635 3965 11640 3985
rect 11660 3965 11665 3985
rect 11635 3960 11665 3965
rect 11640 3955 11660 3960
rect 11550 3870 11570 3875
rect 11545 3865 11575 3870
rect 11545 3845 11550 3865
rect 11570 3845 11575 3865
rect 11545 3840 11575 3845
rect 11505 3830 11525 3835
rect 11500 3825 11530 3830
rect 11500 3805 11505 3825
rect 11525 3805 11530 3825
rect 11500 3800 11530 3805
rect 11005 3620 11035 3625
rect 11005 3600 11010 3620
rect 11030 3600 11035 3620
rect 11005 3595 11035 3600
rect 11185 3620 11215 3625
rect 11185 3600 11190 3620
rect 11210 3600 11215 3620
rect 11185 3595 11215 3600
rect 11365 3620 11395 3625
rect 11365 3600 11370 3620
rect 11390 3600 11395 3620
rect 11365 3595 11395 3600
rect 11010 3590 11030 3595
rect 11190 3590 11210 3595
rect 11370 3590 11390 3595
rect 11505 3575 11525 3800
rect 11550 3625 11570 3840
rect 11545 3620 11575 3625
rect 11545 3600 11550 3620
rect 11570 3600 11575 3620
rect 11545 3595 11575 3600
rect 11550 3590 11570 3595
rect 11685 3575 11705 4080
rect 11820 3990 11840 4165
rect 11910 4110 11930 4115
rect 11905 4105 11935 4110
rect 11905 4085 11910 4105
rect 11930 4085 11935 4105
rect 11905 4080 11935 4085
rect 11815 3985 11845 3990
rect 11815 3965 11820 3985
rect 11840 3965 11845 3985
rect 11815 3960 11845 3965
rect 11820 3955 11840 3960
rect 11730 3870 11750 3875
rect 11725 3865 11755 3870
rect 11725 3845 11730 3865
rect 11750 3845 11755 3865
rect 11725 3840 11755 3845
rect 11730 3625 11750 3840
rect 11865 3830 11885 3835
rect 11860 3825 11890 3830
rect 11860 3805 11865 3825
rect 11885 3805 11890 3825
rect 11860 3800 11890 3805
rect 11725 3620 11755 3625
rect 11725 3600 11730 3620
rect 11750 3600 11755 3620
rect 11725 3595 11755 3600
rect 11730 3590 11750 3595
rect 11865 3575 11885 3800
rect 11910 3625 11930 4080
rect 12000 4030 12020 4165
rect 12090 4110 12110 4115
rect 12085 4105 12115 4110
rect 12085 4085 12090 4105
rect 12110 4085 12115 4105
rect 12085 4080 12115 4085
rect 11995 4025 12025 4030
rect 11995 4005 12000 4025
rect 12020 4005 12025 4025
rect 11995 4000 12025 4005
rect 12000 3995 12020 4000
rect 12045 3830 12065 3835
rect 12040 3825 12070 3830
rect 12040 3805 12045 3825
rect 12065 3805 12070 3825
rect 12040 3800 12070 3805
rect 11905 3620 11935 3625
rect 11905 3600 11910 3620
rect 11930 3600 11935 3620
rect 11905 3595 11935 3600
rect 11910 3590 11930 3595
rect 12045 3575 12065 3800
rect 12090 3625 12110 4080
rect 12180 3790 12200 4165
rect 12225 3950 12245 4215
rect 12360 4195 12380 4200
rect 12355 4190 12385 4195
rect 12355 4170 12360 4190
rect 12380 4170 12385 4190
rect 12355 4165 12385 4170
rect 12220 3945 12250 3950
rect 12220 3925 12225 3945
rect 12245 3925 12250 3945
rect 12220 3920 12250 3925
rect 12225 3915 12245 3920
rect 12270 3910 12290 3915
rect 12360 3910 12380 4165
rect 12405 3910 12425 4215
rect 12540 4195 12560 4200
rect 12535 4190 12565 4195
rect 12535 4170 12540 4190
rect 12560 4170 12565 4190
rect 12535 4165 12565 4170
rect 12450 3910 12470 3915
rect 12540 3910 12560 4165
rect 12585 3950 12605 4215
rect 13305 4210 13325 4215
rect 12720 4195 12740 4200
rect 12900 4195 12920 4200
rect 13080 4195 13100 4200
rect 13260 4195 13280 4200
rect 13440 4195 13460 4200
rect 12715 4190 12745 4195
rect 12715 4170 12720 4190
rect 12740 4170 12745 4190
rect 12715 4165 12745 4170
rect 12895 4190 12925 4195
rect 12895 4170 12900 4190
rect 12920 4170 12925 4190
rect 12895 4165 12925 4170
rect 13075 4190 13105 4195
rect 13075 4170 13080 4190
rect 13100 4170 13105 4190
rect 13075 4165 13105 4170
rect 13255 4190 13285 4195
rect 13255 4170 13260 4190
rect 13280 4170 13285 4190
rect 13255 4165 13285 4170
rect 13435 4190 13465 4195
rect 13435 4170 13440 4190
rect 13460 4170 13465 4190
rect 13435 4165 13465 4170
rect 12630 4110 12650 4115
rect 12625 4105 12655 4110
rect 12625 4085 12630 4105
rect 12650 4085 12655 4105
rect 12625 4080 12655 4085
rect 12580 3945 12610 3950
rect 12580 3925 12585 3945
rect 12605 3925 12610 3945
rect 12580 3920 12610 3925
rect 12585 3915 12605 3920
rect 12265 3905 12295 3910
rect 12265 3885 12270 3905
rect 12290 3885 12295 3905
rect 12265 3880 12295 3885
rect 12355 3905 12385 3910
rect 12355 3885 12360 3905
rect 12380 3885 12385 3905
rect 12355 3880 12385 3885
rect 12400 3905 12430 3910
rect 12400 3885 12405 3905
rect 12425 3885 12430 3905
rect 12400 3880 12430 3885
rect 12445 3905 12475 3910
rect 12445 3885 12450 3905
rect 12470 3885 12475 3905
rect 12445 3880 12475 3885
rect 12535 3905 12565 3910
rect 12535 3885 12540 3905
rect 12560 3885 12565 3905
rect 12535 3880 12565 3885
rect 12175 3785 12205 3790
rect 12175 3765 12180 3785
rect 12200 3765 12205 3785
rect 12175 3760 12205 3765
rect 12180 3755 12200 3760
rect 12270 3625 12290 3880
rect 12360 3875 12380 3880
rect 12085 3620 12115 3625
rect 12085 3600 12090 3620
rect 12110 3600 12115 3620
rect 12085 3595 12115 3600
rect 12265 3620 12295 3625
rect 12265 3600 12270 3620
rect 12290 3600 12295 3620
rect 12265 3595 12295 3600
rect 12090 3590 12110 3595
rect 12270 3590 12290 3595
rect 12405 3575 12425 3880
rect 12450 3625 12470 3880
rect 12540 3875 12560 3880
rect 12630 3625 12650 4080
rect 12720 3790 12740 4165
rect 12900 4160 12920 4165
rect 13080 4160 13100 4165
rect 13260 4160 13280 4165
rect 13440 4160 13460 4165
rect 13485 4160 13505 4215
rect 13620 4195 13640 4200
rect 13800 4195 13820 4200
rect 13980 4195 14000 4200
rect 14160 4195 14180 4200
rect 13615 4190 13645 4195
rect 13615 4170 13620 4190
rect 13640 4170 13645 4190
rect 13615 4165 13645 4170
rect 13795 4190 13825 4195
rect 13795 4170 13800 4190
rect 13820 4170 13825 4190
rect 13795 4165 13825 4170
rect 13975 4190 14005 4195
rect 13975 4170 13980 4190
rect 14000 4170 14005 4190
rect 13975 4165 14005 4170
rect 14155 4190 14185 4195
rect 14155 4170 14160 4190
rect 14180 4170 14185 4190
rect 14155 4165 14185 4170
rect 13620 4160 13640 4165
rect 13800 4160 13820 4165
rect 13980 4160 14000 4165
rect 14160 4160 14180 4165
rect 14205 4160 14225 4215
rect 15465 4210 15485 4215
rect 14340 4195 14360 4200
rect 14520 4195 14540 4200
rect 14700 4195 14720 4200
rect 14880 4195 14900 4200
rect 15060 4195 15080 4200
rect 15240 4195 15260 4200
rect 15420 4195 15440 4200
rect 15600 4195 15620 4200
rect 14335 4190 14365 4195
rect 14335 4170 14340 4190
rect 14360 4170 14365 4190
rect 14335 4165 14365 4170
rect 14515 4190 14545 4195
rect 14515 4170 14520 4190
rect 14540 4170 14545 4190
rect 14515 4165 14545 4170
rect 14695 4190 14725 4195
rect 14695 4170 14700 4190
rect 14720 4170 14725 4190
rect 14695 4165 14725 4170
rect 14875 4190 14905 4195
rect 14875 4170 14880 4190
rect 14900 4170 14905 4190
rect 14875 4165 14905 4170
rect 15055 4190 15085 4195
rect 15055 4170 15060 4190
rect 15080 4170 15085 4190
rect 15055 4165 15085 4170
rect 15235 4190 15265 4195
rect 15235 4170 15240 4190
rect 15260 4170 15265 4190
rect 15235 4165 15265 4170
rect 15415 4190 15445 4195
rect 15415 4170 15420 4190
rect 15440 4170 15445 4190
rect 15415 4165 15445 4170
rect 15595 4190 15625 4195
rect 15595 4170 15600 4190
rect 15620 4170 15625 4190
rect 15595 4165 15625 4170
rect 14340 4160 14360 4165
rect 14520 4160 14540 4165
rect 14700 4160 14720 4165
rect 14880 4160 14900 4165
rect 15060 4160 15080 4165
rect 15240 4160 15260 4165
rect 15420 4160 15440 4165
rect 15600 4160 15620 4165
rect 15645 4160 15665 4215
rect 15780 4195 15800 4200
rect 15960 4195 15980 4200
rect 15775 4190 15805 4195
rect 15775 4170 15780 4190
rect 15800 4170 15805 4190
rect 15775 4165 15805 4170
rect 15955 4190 15985 4195
rect 15955 4170 15960 4190
rect 15980 4170 15985 4190
rect 15955 4165 15985 4170
rect 15780 4160 15800 4165
rect 15960 4160 15980 4165
rect 16005 4160 16025 4215
rect 16140 4195 16160 4200
rect 16320 4195 16340 4200
rect 16135 4190 16165 4195
rect 16135 4170 16140 4190
rect 16160 4170 16165 4190
rect 16135 4165 16165 4170
rect 16315 4190 16345 4195
rect 16315 4170 16320 4190
rect 16340 4170 16345 4190
rect 16315 4165 16345 4170
rect 16140 4160 16160 4165
rect 16320 4160 16340 4165
rect 16365 4160 16385 4215
rect 17625 4210 17645 4215
rect 16500 4195 16520 4200
rect 16680 4195 16700 4200
rect 16860 4195 16880 4200
rect 17040 4195 17060 4200
rect 17220 4195 17240 4200
rect 17400 4195 17420 4200
rect 17580 4195 17600 4200
rect 17760 4195 17780 4200
rect 16495 4190 16525 4195
rect 16495 4170 16500 4190
rect 16520 4170 16525 4190
rect 16495 4165 16525 4170
rect 16675 4190 16705 4195
rect 16675 4170 16680 4190
rect 16700 4170 16705 4190
rect 16675 4165 16705 4170
rect 16855 4190 16885 4195
rect 16855 4170 16860 4190
rect 16880 4170 16885 4190
rect 16855 4165 16885 4170
rect 17035 4190 17065 4195
rect 17035 4170 17040 4190
rect 17060 4170 17065 4190
rect 17035 4165 17065 4170
rect 17215 4190 17245 4195
rect 17215 4170 17220 4190
rect 17240 4170 17245 4190
rect 17215 4165 17245 4170
rect 17395 4190 17425 4195
rect 17395 4170 17400 4190
rect 17420 4170 17425 4190
rect 17395 4165 17425 4170
rect 17575 4190 17605 4195
rect 17575 4170 17580 4190
rect 17600 4170 17605 4190
rect 17575 4165 17605 4170
rect 17755 4190 17785 4195
rect 17755 4170 17760 4190
rect 17780 4170 17785 4190
rect 17755 4165 17785 4170
rect 16500 4160 16520 4165
rect 16680 4160 16700 4165
rect 16860 4160 16880 4165
rect 17040 4160 17060 4165
rect 17220 4160 17240 4165
rect 17400 4160 17420 4165
rect 17580 4160 17600 4165
rect 17760 4160 17780 4165
rect 17805 4160 17825 4215
rect 17940 4195 17960 4200
rect 18120 4195 18140 4200
rect 17935 4190 17965 4195
rect 17935 4170 17940 4190
rect 17960 4170 17965 4190
rect 17935 4165 17965 4170
rect 18115 4190 18145 4195
rect 18115 4170 18120 4190
rect 18140 4170 18145 4190
rect 18115 4165 18145 4170
rect 17940 4160 17960 4165
rect 18120 4160 18140 4165
rect 18165 4160 18185 4215
rect 18300 4195 18320 4200
rect 18480 4195 18500 4200
rect 18295 4190 18325 4195
rect 18295 4170 18300 4190
rect 18320 4170 18325 4190
rect 18295 4165 18325 4170
rect 18475 4190 18505 4195
rect 18475 4170 18480 4190
rect 18500 4170 18505 4190
rect 18475 4165 18505 4170
rect 18300 4160 18320 4165
rect 18480 4160 18500 4165
rect 18525 4160 18545 4215
rect 18660 4195 18680 4200
rect 18840 4195 18860 4200
rect 19020 4195 19040 4200
rect 19200 4195 19220 4200
rect 18655 4190 18685 4195
rect 18655 4170 18660 4190
rect 18680 4170 18685 4190
rect 18655 4165 18685 4170
rect 18835 4190 18865 4195
rect 18835 4170 18840 4190
rect 18860 4170 18865 4190
rect 18835 4165 18865 4170
rect 19015 4190 19045 4195
rect 19015 4170 19020 4190
rect 19040 4170 19045 4190
rect 19015 4165 19045 4170
rect 19195 4190 19225 4195
rect 19195 4170 19200 4190
rect 19220 4170 19225 4190
rect 19195 4165 19225 4170
rect 18660 4160 18680 4165
rect 18840 4160 18860 4165
rect 19020 4160 19040 4165
rect 19200 4160 19220 4165
rect 19335 4160 19355 4215
rect 19380 4195 19400 4200
rect 19375 4190 19405 4195
rect 19375 4170 19380 4190
rect 19400 4170 19405 4190
rect 19375 4165 19405 4170
rect 19380 4160 19400 4165
rect 19515 4160 19535 4215
rect 19560 4195 19580 4200
rect 19555 4190 19585 4195
rect 19555 4170 19560 4190
rect 19580 4170 19585 4190
rect 19555 4165 19585 4170
rect 19560 4160 19580 4165
rect 19695 4160 19715 4215
rect 19740 4195 19760 4200
rect 19735 4190 19765 4195
rect 19735 4170 19740 4190
rect 19760 4170 19765 4190
rect 19735 4165 19765 4170
rect 19740 4160 19760 4165
rect 19875 4160 19895 4215
rect 19920 4195 19940 4200
rect 19915 4190 19945 4195
rect 19915 4170 19920 4190
rect 19940 4170 19945 4190
rect 19915 4165 19945 4170
rect 19920 4160 19940 4165
rect 20055 4075 20075 4215
rect 20145 4110 20165 4215
rect 20140 4105 20170 4110
rect 20140 4085 20145 4105
rect 20165 4085 20170 4105
rect 20140 4080 20170 4085
rect 20145 4075 20165 4080
rect 20235 3910 20255 4215
rect 20325 3990 20345 4215
rect 20320 3985 20350 3990
rect 20320 3965 20325 3985
rect 20345 3965 20350 3985
rect 20320 3960 20350 3965
rect 20230 3905 20260 3910
rect 20230 3885 20235 3905
rect 20255 3885 20260 3905
rect 20230 3880 20260 3885
rect 12715 3785 12745 3790
rect 12715 3765 12720 3785
rect 12740 3765 12745 3785
rect 12715 3760 12745 3765
rect 12720 3755 12740 3760
rect 12810 3625 12830 3630
rect 12990 3625 13010 3630
rect 13170 3625 13190 3630
rect 13350 3625 13370 3630
rect 12445 3620 12475 3625
rect 12445 3600 12450 3620
rect 12470 3600 12475 3620
rect 12445 3595 12475 3600
rect 12625 3620 12655 3625
rect 12625 3600 12630 3620
rect 12650 3600 12655 3620
rect 12625 3595 12655 3600
rect 12805 3620 12835 3625
rect 12805 3600 12810 3620
rect 12830 3600 12835 3620
rect 12805 3595 12835 3600
rect 12985 3620 13015 3625
rect 12985 3600 12990 3620
rect 13010 3600 13015 3620
rect 12985 3595 13015 3600
rect 13165 3620 13195 3625
rect 13165 3600 13170 3620
rect 13190 3600 13195 3620
rect 13165 3595 13195 3600
rect 13345 3620 13375 3625
rect 13345 3600 13350 3620
rect 13370 3600 13375 3620
rect 13345 3595 13375 3600
rect 12450 3590 12470 3595
rect 12630 3590 12650 3595
rect 12810 3590 12830 3595
rect 12990 3590 13010 3595
rect 13170 3590 13190 3595
rect 13350 3590 13370 3595
rect 13485 3575 13505 3630
rect 13530 3625 13550 3630
rect 13710 3625 13730 3630
rect 13525 3620 13555 3625
rect 13525 3600 13530 3620
rect 13550 3600 13555 3620
rect 13525 3595 13555 3600
rect 13705 3620 13735 3625
rect 13705 3600 13710 3620
rect 13730 3600 13735 3620
rect 13705 3595 13735 3600
rect 13530 3590 13550 3595
rect 13710 3590 13730 3595
rect 13845 3575 13865 3630
rect 13890 3625 13910 3630
rect 14070 3625 14090 3630
rect 13885 3620 13915 3625
rect 13885 3600 13890 3620
rect 13910 3600 13915 3620
rect 13885 3595 13915 3600
rect 14065 3620 14095 3625
rect 14065 3600 14070 3620
rect 14090 3600 14095 3620
rect 14065 3595 14095 3600
rect 13890 3590 13910 3595
rect 14070 3590 14090 3595
rect 14205 3575 14225 3630
rect 14250 3625 14270 3630
rect 14430 3625 14450 3630
rect 14610 3625 14630 3630
rect 14790 3625 14810 3630
rect 14970 3625 14990 3630
rect 15150 3625 15170 3630
rect 15330 3625 15350 3630
rect 15510 3625 15530 3630
rect 14245 3620 14275 3625
rect 14245 3600 14250 3620
rect 14270 3600 14275 3620
rect 14245 3595 14275 3600
rect 14425 3620 14455 3625
rect 14425 3600 14430 3620
rect 14450 3600 14455 3620
rect 14425 3595 14455 3600
rect 14605 3620 14635 3625
rect 14605 3600 14610 3620
rect 14630 3600 14635 3620
rect 14605 3595 14635 3600
rect 14785 3620 14815 3625
rect 14785 3600 14790 3620
rect 14810 3600 14815 3620
rect 14785 3595 14815 3600
rect 14965 3620 14995 3625
rect 14965 3600 14970 3620
rect 14990 3600 14995 3620
rect 14965 3595 14995 3600
rect 15145 3620 15175 3625
rect 15145 3600 15150 3620
rect 15170 3600 15175 3620
rect 15145 3595 15175 3600
rect 15325 3620 15355 3625
rect 15325 3600 15330 3620
rect 15350 3600 15355 3620
rect 15325 3595 15355 3600
rect 15505 3620 15535 3625
rect 15505 3600 15510 3620
rect 15530 3600 15535 3620
rect 15505 3595 15535 3600
rect 14250 3590 14270 3595
rect 14430 3590 14450 3595
rect 14610 3590 14630 3595
rect 14790 3590 14810 3595
rect 14970 3590 14990 3595
rect 15150 3590 15170 3595
rect 15330 3590 15350 3595
rect 15510 3590 15530 3595
rect 15645 3575 15665 3630
rect 15690 3625 15710 3630
rect 15870 3625 15890 3630
rect 16050 3625 16070 3630
rect 16230 3625 16250 3630
rect 15685 3620 15715 3625
rect 15685 3600 15690 3620
rect 15710 3600 15715 3620
rect 15685 3595 15715 3600
rect 15865 3620 15895 3625
rect 15865 3600 15870 3620
rect 15890 3600 15895 3620
rect 15865 3595 15895 3600
rect 16045 3620 16075 3625
rect 16045 3600 16050 3620
rect 16070 3600 16075 3620
rect 16045 3595 16075 3600
rect 16225 3620 16255 3625
rect 16225 3600 16230 3620
rect 16250 3600 16255 3620
rect 16225 3595 16255 3600
rect 15690 3590 15710 3595
rect 15870 3590 15890 3595
rect 16050 3590 16070 3595
rect 16230 3590 16250 3595
rect 16365 3575 16385 3630
rect 16410 3625 16430 3630
rect 16590 3625 16610 3630
rect 16770 3625 16790 3630
rect 16950 3625 16970 3630
rect 17130 3625 17150 3630
rect 17310 3625 17330 3630
rect 17490 3625 17510 3630
rect 17670 3625 17690 3630
rect 16405 3620 16435 3625
rect 16405 3600 16410 3620
rect 16430 3600 16435 3620
rect 16405 3595 16435 3600
rect 16585 3620 16615 3625
rect 16585 3600 16590 3620
rect 16610 3600 16615 3620
rect 16585 3595 16615 3600
rect 16765 3620 16795 3625
rect 16765 3600 16770 3620
rect 16790 3600 16795 3620
rect 16765 3595 16795 3600
rect 16945 3620 16975 3625
rect 16945 3600 16950 3620
rect 16970 3600 16975 3620
rect 16945 3595 16975 3600
rect 17125 3620 17155 3625
rect 17125 3600 17130 3620
rect 17150 3600 17155 3620
rect 17125 3595 17155 3600
rect 17305 3620 17335 3625
rect 17305 3600 17310 3620
rect 17330 3600 17335 3620
rect 17305 3595 17335 3600
rect 17485 3620 17515 3625
rect 17485 3600 17490 3620
rect 17510 3600 17515 3620
rect 17485 3595 17515 3600
rect 17665 3620 17695 3625
rect 17665 3600 17670 3620
rect 17690 3600 17695 3620
rect 17665 3595 17695 3600
rect 16410 3590 16430 3595
rect 16590 3590 16610 3595
rect 16770 3590 16790 3595
rect 16950 3590 16970 3595
rect 17130 3590 17150 3595
rect 17310 3590 17330 3595
rect 17490 3590 17510 3595
rect 17670 3590 17690 3595
rect 17805 3575 17825 3630
rect 17850 3625 17870 3630
rect 18030 3625 18050 3630
rect 18210 3625 18230 3630
rect 18390 3625 18410 3630
rect 17845 3620 17875 3625
rect 17845 3600 17850 3620
rect 17870 3600 17875 3620
rect 17845 3595 17875 3600
rect 18025 3620 18055 3625
rect 18025 3600 18030 3620
rect 18050 3600 18055 3620
rect 18025 3595 18055 3600
rect 18205 3620 18235 3625
rect 18205 3600 18210 3620
rect 18230 3600 18235 3620
rect 18205 3595 18235 3600
rect 18385 3620 18415 3625
rect 18385 3600 18390 3620
rect 18410 3600 18415 3620
rect 18385 3595 18415 3600
rect 17850 3590 17870 3595
rect 18030 3590 18050 3595
rect 18210 3590 18230 3595
rect 18390 3590 18410 3595
rect 18525 3575 18545 3630
rect 18570 3625 18590 3630
rect 18750 3625 18770 3630
rect 18930 3625 18950 3630
rect 19110 3625 19130 3630
rect 19290 3625 19310 3630
rect 18565 3620 18595 3625
rect 18565 3600 18570 3620
rect 18590 3600 18595 3620
rect 18565 3595 18595 3600
rect 18745 3620 18775 3625
rect 18745 3600 18750 3620
rect 18770 3600 18775 3620
rect 18745 3595 18775 3600
rect 18925 3620 18955 3625
rect 18925 3600 18930 3620
rect 18950 3600 18955 3620
rect 18925 3595 18955 3600
rect 19105 3620 19135 3625
rect 19105 3600 19110 3620
rect 19130 3600 19135 3620
rect 19105 3595 19135 3600
rect 19285 3620 19315 3625
rect 19285 3600 19290 3620
rect 19310 3600 19315 3620
rect 19285 3595 19315 3600
rect 18570 3590 18590 3595
rect 18750 3590 18770 3595
rect 18930 3590 18950 3595
rect 19110 3590 19130 3595
rect 19290 3590 19310 3595
rect 19335 3575 19355 3630
rect 19470 3625 19490 3630
rect 19465 3620 19495 3625
rect 19465 3600 19470 3620
rect 19490 3600 19495 3620
rect 19465 3595 19495 3600
rect 19470 3590 19490 3595
rect 19515 3575 19535 3630
rect 19650 3625 19670 3630
rect 19645 3620 19675 3625
rect 19645 3600 19650 3620
rect 19670 3600 19675 3620
rect 19645 3595 19675 3600
rect 19650 3590 19670 3595
rect 19695 3575 19715 3630
rect 19830 3625 19850 3630
rect 19825 3620 19855 3625
rect 19825 3600 19830 3620
rect 19850 3600 19855 3620
rect 19825 3595 19855 3600
rect 19830 3590 19850 3595
rect 19875 3575 19895 3630
rect 20055 3575 20075 3630
rect 20145 3575 20165 3630
rect 20235 3575 20255 3880
rect 20325 3575 20345 3960
rect 20415 3950 20435 4215
rect 20410 3945 20440 3950
rect 20410 3925 20415 3945
rect 20435 3925 20440 3945
rect 20410 3920 20440 3925
rect 20415 3575 20435 3920
rect 20505 3750 20525 4215
rect 20500 3745 20530 3750
rect 20500 3725 20505 3745
rect 20525 3725 20530 3745
rect 20500 3720 20530 3725
rect 20505 3575 20525 3720
rect 20595 3710 20615 4215
rect 20590 3705 20620 3710
rect 20590 3685 20595 3705
rect 20615 3685 20620 3705
rect 20590 3680 20620 3685
rect 20595 3575 20615 3680
rect 9160 3565 9190 3575
rect 9160 3485 9165 3565
rect 9185 3485 9190 3565
rect 9160 3475 9190 3485
rect 9250 3475 9280 3575
rect 9340 3475 9370 3575
rect 9430 3475 9460 3575
rect 9520 3475 9550 3575
rect 9610 3475 9640 3575
rect 9700 3475 9730 3575
rect 9790 3475 9820 3575
rect 9880 3565 9910 3575
rect 9880 3485 9885 3565
rect 9905 3485 9910 3565
rect 9880 3475 9910 3485
rect 9970 3565 10000 3575
rect 9970 3485 9975 3565
rect 9995 3485 10000 3565
rect 9970 3475 10000 3485
rect 10060 3565 10090 3575
rect 10060 3485 10065 3565
rect 10085 3485 10090 3565
rect 10060 3475 10090 3485
rect 10150 3565 10180 3575
rect 10150 3485 10155 3565
rect 10175 3485 10180 3565
rect 10150 3475 10180 3485
rect 10240 3565 10270 3575
rect 10240 3485 10245 3565
rect 10265 3485 10270 3565
rect 10240 3475 10270 3485
rect 10330 3565 10360 3575
rect 10330 3485 10335 3565
rect 10355 3485 10360 3565
rect 10330 3475 10360 3485
rect 10420 3565 10450 3575
rect 10420 3485 10425 3565
rect 10445 3485 10450 3565
rect 10420 3475 10450 3485
rect 10510 3565 10540 3575
rect 10510 3485 10515 3565
rect 10535 3485 10540 3565
rect 10510 3475 10540 3485
rect 10600 3565 10630 3575
rect 10600 3485 10605 3565
rect 10625 3485 10630 3565
rect 10600 3475 10630 3485
rect 10690 3565 10720 3575
rect 10690 3485 10695 3565
rect 10715 3485 10720 3565
rect 10690 3475 10720 3485
rect 10780 3565 10810 3575
rect 10780 3485 10785 3565
rect 10805 3485 10810 3565
rect 10780 3475 10810 3485
rect 10870 3565 10900 3575
rect 10870 3485 10875 3565
rect 10895 3485 10900 3565
rect 10870 3475 10900 3485
rect 10960 3565 10990 3575
rect 10960 3485 10965 3565
rect 10985 3485 10990 3565
rect 10960 3475 10990 3485
rect 11050 3565 11080 3575
rect 11050 3485 11055 3565
rect 11075 3485 11080 3565
rect 11050 3475 11080 3485
rect 11140 3565 11170 3575
rect 11140 3485 11145 3565
rect 11165 3485 11170 3565
rect 11140 3475 11170 3485
rect 11230 3565 11260 3575
rect 11230 3485 11235 3565
rect 11255 3485 11260 3565
rect 11230 3475 11260 3485
rect 11320 3565 11350 3575
rect 11320 3485 11325 3565
rect 11345 3485 11350 3565
rect 11320 3475 11350 3485
rect 11410 3565 11440 3575
rect 11410 3485 11415 3565
rect 11435 3485 11440 3565
rect 11410 3475 11440 3485
rect 11500 3565 11530 3575
rect 11500 3485 11505 3565
rect 11525 3485 11530 3565
rect 11500 3475 11530 3485
rect 11590 3565 11620 3575
rect 11590 3485 11595 3565
rect 11615 3485 11620 3565
rect 11590 3475 11620 3485
rect 11680 3565 11710 3575
rect 11680 3485 11685 3565
rect 11705 3485 11710 3565
rect 11680 3475 11710 3485
rect 11770 3565 11800 3575
rect 11770 3485 11775 3565
rect 11795 3485 11800 3565
rect 11770 3475 11800 3485
rect 11860 3565 11890 3575
rect 11860 3485 11865 3565
rect 11885 3485 11890 3565
rect 11860 3475 11890 3485
rect 11950 3565 11980 3575
rect 11950 3485 11955 3565
rect 11975 3485 11980 3565
rect 11950 3475 11980 3485
rect 12040 3565 12070 3575
rect 12040 3485 12045 3565
rect 12065 3485 12070 3565
rect 12040 3475 12070 3485
rect 12130 3565 12160 3575
rect 12130 3485 12135 3565
rect 12155 3485 12160 3565
rect 12130 3475 12160 3485
rect 12220 3565 12250 3575
rect 12220 3485 12225 3565
rect 12245 3485 12250 3565
rect 12220 3475 12250 3485
rect 12310 3565 12340 3575
rect 12310 3485 12315 3565
rect 12335 3485 12340 3565
rect 12310 3475 12340 3485
rect 12400 3565 12430 3575
rect 12400 3485 12405 3565
rect 12425 3485 12430 3565
rect 12400 3475 12430 3485
rect 12490 3565 12520 3575
rect 12490 3485 12495 3565
rect 12515 3485 12520 3565
rect 12490 3475 12520 3485
rect 12580 3565 12610 3575
rect 12580 3485 12585 3565
rect 12605 3485 12610 3565
rect 12580 3475 12610 3485
rect 12670 3565 12700 3575
rect 12670 3485 12675 3565
rect 12695 3485 12700 3565
rect 12670 3475 12700 3485
rect 12760 3565 12790 3575
rect 12760 3485 12765 3565
rect 12785 3485 12790 3565
rect 12760 3475 12790 3485
rect 12850 3565 12880 3575
rect 12850 3485 12855 3565
rect 12875 3485 12880 3565
rect 12850 3475 12880 3485
rect 12940 3565 12970 3575
rect 12940 3485 12945 3565
rect 12965 3485 12970 3565
rect 12940 3475 12970 3485
rect 13030 3565 13060 3575
rect 13030 3485 13035 3565
rect 13055 3485 13060 3565
rect 13030 3475 13060 3485
rect 13120 3565 13150 3575
rect 13120 3485 13125 3565
rect 13145 3485 13150 3565
rect 13120 3475 13150 3485
rect 13210 3565 13240 3575
rect 13210 3485 13215 3565
rect 13235 3485 13240 3565
rect 13210 3475 13240 3485
rect 13300 3565 13330 3575
rect 13300 3485 13305 3565
rect 13325 3485 13330 3565
rect 13300 3475 13330 3485
rect 13390 3565 13420 3575
rect 13390 3485 13395 3565
rect 13415 3485 13420 3565
rect 13390 3475 13420 3485
rect 13480 3565 13510 3575
rect 13480 3485 13485 3565
rect 13505 3485 13510 3565
rect 13480 3475 13510 3485
rect 13570 3565 13600 3575
rect 13570 3485 13575 3565
rect 13595 3485 13600 3565
rect 13570 3475 13600 3485
rect 13660 3565 13690 3575
rect 13660 3485 13665 3565
rect 13685 3485 13690 3565
rect 13660 3475 13690 3485
rect 13750 3565 13780 3575
rect 13750 3485 13755 3565
rect 13775 3485 13780 3565
rect 13750 3475 13780 3485
rect 13840 3565 13870 3575
rect 13840 3485 13845 3565
rect 13865 3485 13870 3565
rect 13840 3475 13870 3485
rect 13930 3565 13960 3575
rect 13930 3485 13935 3565
rect 13955 3485 13960 3565
rect 13930 3475 13960 3485
rect 14020 3565 14050 3575
rect 14020 3485 14025 3565
rect 14045 3485 14050 3565
rect 14020 3475 14050 3485
rect 14110 3565 14140 3575
rect 14110 3485 14115 3565
rect 14135 3485 14140 3565
rect 14110 3475 14140 3485
rect 14200 3565 14230 3575
rect 14200 3485 14205 3565
rect 14225 3485 14230 3565
rect 14200 3475 14230 3485
rect 14290 3565 14320 3575
rect 14290 3485 14295 3565
rect 14315 3485 14320 3565
rect 14290 3475 14320 3485
rect 14380 3565 14410 3575
rect 14380 3485 14385 3565
rect 14405 3485 14410 3565
rect 14380 3475 14410 3485
rect 14470 3565 14500 3575
rect 14470 3485 14475 3565
rect 14495 3485 14500 3565
rect 14470 3475 14500 3485
rect 14560 3565 14590 3575
rect 14560 3485 14565 3565
rect 14585 3485 14590 3565
rect 14560 3475 14590 3485
rect 14650 3565 14680 3575
rect 14650 3485 14655 3565
rect 14675 3485 14680 3565
rect 14650 3475 14680 3485
rect 14740 3565 14770 3575
rect 14740 3485 14745 3565
rect 14765 3485 14770 3565
rect 14740 3475 14770 3485
rect 14830 3565 14860 3575
rect 14830 3485 14835 3565
rect 14855 3485 14860 3565
rect 14830 3475 14860 3485
rect 14920 3565 14950 3575
rect 14920 3485 14925 3565
rect 14945 3485 14950 3565
rect 14920 3475 14950 3485
rect 15010 3565 15040 3575
rect 15010 3485 15015 3565
rect 15035 3485 15040 3565
rect 15010 3475 15040 3485
rect 15100 3565 15130 3575
rect 15100 3485 15105 3565
rect 15125 3485 15130 3565
rect 15100 3475 15130 3485
rect 15190 3565 15220 3575
rect 15190 3485 15195 3565
rect 15215 3485 15220 3565
rect 15190 3475 15220 3485
rect 15280 3565 15310 3575
rect 15280 3485 15285 3565
rect 15305 3485 15310 3565
rect 15280 3475 15310 3485
rect 15370 3565 15400 3575
rect 15370 3485 15375 3565
rect 15395 3485 15400 3565
rect 15370 3475 15400 3485
rect 15460 3565 15490 3575
rect 15460 3485 15465 3565
rect 15485 3485 15490 3565
rect 15460 3475 15490 3485
rect 15550 3565 15580 3575
rect 15550 3485 15555 3565
rect 15575 3485 15580 3565
rect 15550 3475 15580 3485
rect 15640 3565 15670 3575
rect 15640 3485 15645 3565
rect 15665 3485 15670 3565
rect 15640 3475 15670 3485
rect 15730 3565 15760 3575
rect 15730 3485 15735 3565
rect 15755 3485 15760 3565
rect 15730 3475 15760 3485
rect 15820 3565 15850 3575
rect 15820 3485 15825 3565
rect 15845 3485 15850 3565
rect 15820 3475 15850 3485
rect 15910 3565 15940 3575
rect 15910 3485 15915 3565
rect 15935 3485 15940 3565
rect 15910 3475 15940 3485
rect 16000 3565 16030 3575
rect 16000 3485 16005 3565
rect 16025 3485 16030 3565
rect 16000 3475 16030 3485
rect 16090 3565 16120 3575
rect 16090 3485 16095 3565
rect 16115 3485 16120 3565
rect 16090 3475 16120 3485
rect 16180 3565 16210 3575
rect 16180 3485 16185 3565
rect 16205 3485 16210 3565
rect 16180 3475 16210 3485
rect 16270 3565 16300 3575
rect 16270 3485 16275 3565
rect 16295 3485 16300 3565
rect 16270 3475 16300 3485
rect 16360 3565 16390 3575
rect 16360 3485 16365 3565
rect 16385 3485 16390 3565
rect 16360 3475 16390 3485
rect 16450 3565 16480 3575
rect 16450 3485 16455 3565
rect 16475 3485 16480 3565
rect 16450 3475 16480 3485
rect 16540 3565 16570 3575
rect 16540 3485 16545 3565
rect 16565 3485 16570 3565
rect 16540 3475 16570 3485
rect 16630 3565 16660 3575
rect 16630 3485 16635 3565
rect 16655 3485 16660 3565
rect 16630 3475 16660 3485
rect 16720 3565 16750 3575
rect 16720 3485 16725 3565
rect 16745 3485 16750 3565
rect 16720 3475 16750 3485
rect 16810 3565 16840 3575
rect 16810 3485 16815 3565
rect 16835 3485 16840 3565
rect 16810 3475 16840 3485
rect 16900 3565 16930 3575
rect 16900 3485 16905 3565
rect 16925 3485 16930 3565
rect 16900 3475 16930 3485
rect 16990 3565 17020 3575
rect 16990 3485 16995 3565
rect 17015 3485 17020 3565
rect 16990 3475 17020 3485
rect 17080 3565 17110 3575
rect 17080 3485 17085 3565
rect 17105 3485 17110 3565
rect 17080 3475 17110 3485
rect 17170 3565 17200 3575
rect 17170 3485 17175 3565
rect 17195 3485 17200 3565
rect 17170 3475 17200 3485
rect 17260 3565 17290 3575
rect 17260 3485 17265 3565
rect 17285 3485 17290 3565
rect 17260 3475 17290 3485
rect 17350 3565 17380 3575
rect 17350 3485 17355 3565
rect 17375 3485 17380 3565
rect 17350 3475 17380 3485
rect 17440 3565 17470 3575
rect 17440 3485 17445 3565
rect 17465 3485 17470 3565
rect 17440 3475 17470 3485
rect 17530 3565 17560 3575
rect 17530 3485 17535 3565
rect 17555 3485 17560 3565
rect 17530 3475 17560 3485
rect 17620 3565 17650 3575
rect 17620 3485 17625 3565
rect 17645 3485 17650 3565
rect 17620 3475 17650 3485
rect 17710 3565 17740 3575
rect 17710 3485 17715 3565
rect 17735 3485 17740 3565
rect 17710 3475 17740 3485
rect 17800 3565 17830 3575
rect 17800 3485 17805 3565
rect 17825 3485 17830 3565
rect 17800 3475 17830 3485
rect 17890 3565 17920 3575
rect 17890 3485 17895 3565
rect 17915 3485 17920 3565
rect 17890 3475 17920 3485
rect 17980 3565 18010 3575
rect 17980 3485 17985 3565
rect 18005 3485 18010 3565
rect 17980 3475 18010 3485
rect 18070 3565 18100 3575
rect 18070 3485 18075 3565
rect 18095 3485 18100 3565
rect 18070 3475 18100 3485
rect 18160 3565 18190 3575
rect 18160 3485 18165 3565
rect 18185 3485 18190 3565
rect 18160 3475 18190 3485
rect 18250 3565 18280 3575
rect 18250 3485 18255 3565
rect 18275 3485 18280 3565
rect 18250 3475 18280 3485
rect 18340 3565 18370 3575
rect 18340 3485 18345 3565
rect 18365 3485 18370 3565
rect 18340 3475 18370 3485
rect 18430 3565 18460 3575
rect 18430 3485 18435 3565
rect 18455 3485 18460 3565
rect 18430 3475 18460 3485
rect 18520 3565 18550 3575
rect 18520 3485 18525 3565
rect 18545 3485 18550 3565
rect 18520 3475 18550 3485
rect 18610 3565 18640 3575
rect 18610 3485 18615 3565
rect 18635 3485 18640 3565
rect 18610 3475 18640 3485
rect 18700 3565 18730 3575
rect 18700 3485 18705 3565
rect 18725 3485 18730 3565
rect 18700 3475 18730 3485
rect 18790 3565 18820 3575
rect 18790 3485 18795 3565
rect 18815 3485 18820 3565
rect 18790 3475 18820 3485
rect 18880 3565 18910 3575
rect 18880 3485 18885 3565
rect 18905 3485 18910 3565
rect 18880 3475 18910 3485
rect 18970 3565 19000 3575
rect 18970 3485 18975 3565
rect 18995 3485 19000 3565
rect 18970 3475 19000 3485
rect 19060 3565 19090 3575
rect 19060 3485 19065 3565
rect 19085 3485 19090 3565
rect 19060 3475 19090 3485
rect 19150 3565 19180 3575
rect 19150 3485 19155 3565
rect 19175 3485 19180 3565
rect 19150 3475 19180 3485
rect 19240 3565 19270 3575
rect 19240 3485 19245 3565
rect 19265 3485 19270 3565
rect 19240 3475 19270 3485
rect 19330 3565 19360 3575
rect 19330 3485 19335 3565
rect 19355 3485 19360 3565
rect 19330 3475 19360 3485
rect 19420 3565 19450 3575
rect 19420 3485 19425 3565
rect 19445 3485 19450 3565
rect 19420 3475 19450 3485
rect 19510 3565 19540 3575
rect 19510 3485 19515 3565
rect 19535 3485 19540 3565
rect 19510 3475 19540 3485
rect 19600 3565 19630 3575
rect 19600 3485 19605 3565
rect 19625 3485 19630 3565
rect 19600 3475 19630 3485
rect 19690 3565 19720 3575
rect 19690 3485 19695 3565
rect 19715 3485 19720 3565
rect 19690 3475 19720 3485
rect 19780 3565 19810 3575
rect 19780 3485 19785 3565
rect 19805 3485 19810 3565
rect 19780 3475 19810 3485
rect 19870 3565 19900 3575
rect 19870 3485 19875 3565
rect 19895 3485 19900 3565
rect 19870 3475 19900 3485
rect 19960 3565 19990 3575
rect 19960 3485 19965 3565
rect 19985 3485 19990 3565
rect 19960 3475 19990 3485
rect 20050 3475 20080 3575
rect 20140 3475 20170 3575
rect 20230 3475 20260 3575
rect 20320 3475 20350 3575
rect 20410 3475 20440 3575
rect 20500 3475 20530 3575
rect 20590 3475 20620 3575
rect 20680 3565 20710 3575
rect 20680 3485 20685 3565
rect 20705 3485 20710 3565
rect 20680 3475 20710 3485
rect 9165 3455 9185 3475
rect 9885 3455 9905 3475
rect 10605 3455 10625 3475
rect 11325 3455 11345 3475
rect 12045 3455 12065 3475
rect 12765 3455 12785 3475
rect 14925 3455 14945 3475
rect 17085 3455 17105 3475
rect 19245 3455 19265 3475
rect 19425 3455 19445 3475
rect 19605 3455 19625 3475
rect 19785 3455 19805 3475
rect 19965 3455 19985 3475
rect 20685 3455 20705 3475
rect 9020 3420 9025 3450
rect 9055 3420 9060 3450
rect 9020 3415 9060 3420
rect 9155 3450 9195 3455
rect 9155 3420 9160 3450
rect 9190 3420 9195 3450
rect 9155 3415 9195 3420
rect 9875 3450 9915 3455
rect 9875 3420 9880 3450
rect 9910 3420 9915 3450
rect 9875 3415 9915 3420
rect 10055 3450 10095 3455
rect 10055 3420 10060 3450
rect 10090 3420 10095 3450
rect 10055 3415 10095 3420
rect 10235 3450 10275 3455
rect 10235 3420 10240 3450
rect 10270 3420 10275 3450
rect 10235 3415 10275 3420
rect 10415 3450 10455 3455
rect 10415 3420 10420 3450
rect 10450 3420 10455 3450
rect 10415 3415 10455 3420
rect 10595 3450 10635 3455
rect 10595 3420 10600 3450
rect 10630 3420 10635 3450
rect 10595 3415 10635 3420
rect 10775 3450 10815 3455
rect 10775 3420 10780 3450
rect 10810 3420 10815 3450
rect 10775 3415 10815 3420
rect 10955 3450 10995 3455
rect 10955 3420 10960 3450
rect 10990 3420 10995 3450
rect 10955 3415 10995 3420
rect 11135 3450 11175 3455
rect 11135 3420 11140 3450
rect 11170 3420 11175 3450
rect 11135 3415 11175 3420
rect 11315 3450 11355 3455
rect 11315 3420 11320 3450
rect 11350 3420 11355 3450
rect 11315 3415 11355 3420
rect 11495 3450 11535 3455
rect 11495 3420 11500 3450
rect 11530 3420 11535 3450
rect 11495 3415 11535 3420
rect 11675 3450 11715 3455
rect 11675 3420 11680 3450
rect 11710 3420 11715 3450
rect 11675 3415 11715 3420
rect 11855 3450 11895 3455
rect 11855 3420 11860 3450
rect 11890 3420 11895 3450
rect 11855 3415 11895 3420
rect 12035 3450 12075 3455
rect 12035 3420 12040 3450
rect 12070 3420 12075 3450
rect 12035 3415 12075 3420
rect 12215 3450 12255 3455
rect 12215 3420 12220 3450
rect 12250 3420 12255 3450
rect 12215 3415 12255 3420
rect 12395 3450 12435 3455
rect 12395 3420 12400 3450
rect 12430 3420 12435 3450
rect 12395 3415 12435 3420
rect 12575 3450 12615 3455
rect 12575 3420 12580 3450
rect 12610 3420 12615 3450
rect 12575 3415 12615 3420
rect 12755 3450 12795 3455
rect 12755 3420 12760 3450
rect 12790 3420 12795 3450
rect 12755 3415 12795 3420
rect 12935 3450 12975 3455
rect 12935 3420 12940 3450
rect 12970 3420 12975 3450
rect 12935 3415 12975 3420
rect 13115 3450 13155 3455
rect 13115 3420 13120 3450
rect 13150 3420 13155 3450
rect 13115 3415 13155 3420
rect 13295 3450 13335 3455
rect 13295 3420 13300 3450
rect 13330 3420 13335 3450
rect 13295 3415 13335 3420
rect 13475 3450 13515 3455
rect 13475 3420 13480 3450
rect 13510 3420 13515 3450
rect 13475 3415 13515 3420
rect 13655 3450 13695 3455
rect 13655 3420 13660 3450
rect 13690 3420 13695 3450
rect 13655 3415 13695 3420
rect 13835 3450 13875 3455
rect 13835 3420 13840 3450
rect 13870 3420 13875 3450
rect 13835 3415 13875 3420
rect 14015 3450 14055 3455
rect 14015 3420 14020 3450
rect 14050 3420 14055 3450
rect 14015 3415 14055 3420
rect 14195 3450 14235 3455
rect 14195 3420 14200 3450
rect 14230 3420 14235 3450
rect 14195 3415 14235 3420
rect 14375 3450 14415 3455
rect 14375 3420 14380 3450
rect 14410 3420 14415 3450
rect 14375 3415 14415 3420
rect 14555 3450 14595 3455
rect 14555 3420 14560 3450
rect 14590 3420 14595 3450
rect 14555 3415 14595 3420
rect 14735 3450 14775 3455
rect 14735 3420 14740 3450
rect 14770 3420 14775 3450
rect 14735 3415 14775 3420
rect 14915 3450 14955 3455
rect 14915 3420 14920 3450
rect 14950 3420 14955 3450
rect 14915 3415 14955 3420
rect 15095 3450 15135 3455
rect 15095 3420 15100 3450
rect 15130 3420 15135 3450
rect 15095 3415 15135 3420
rect 15275 3450 15315 3455
rect 15275 3420 15280 3450
rect 15310 3420 15315 3450
rect 15275 3415 15315 3420
rect 15455 3450 15495 3455
rect 15455 3420 15460 3450
rect 15490 3420 15495 3450
rect 15455 3415 15495 3420
rect 15635 3450 15675 3455
rect 15635 3420 15640 3450
rect 15670 3420 15675 3450
rect 15635 3415 15675 3420
rect 15815 3450 15855 3455
rect 15815 3420 15820 3450
rect 15850 3420 15855 3450
rect 15815 3415 15855 3420
rect 15995 3450 16035 3455
rect 15995 3420 16000 3450
rect 16030 3420 16035 3450
rect 15995 3415 16035 3420
rect 16175 3450 16215 3455
rect 16175 3420 16180 3450
rect 16210 3420 16215 3450
rect 16175 3415 16215 3420
rect 16355 3450 16395 3455
rect 16355 3420 16360 3450
rect 16390 3420 16395 3450
rect 16355 3415 16395 3420
rect 16535 3450 16575 3455
rect 16535 3420 16540 3450
rect 16570 3420 16575 3450
rect 16535 3415 16575 3420
rect 16715 3450 16755 3455
rect 16715 3420 16720 3450
rect 16750 3420 16755 3450
rect 16715 3415 16755 3420
rect 16895 3450 16935 3455
rect 16895 3420 16900 3450
rect 16930 3420 16935 3450
rect 16895 3415 16935 3420
rect 17075 3450 17115 3455
rect 17075 3420 17080 3450
rect 17110 3420 17115 3450
rect 17075 3415 17115 3420
rect 17255 3450 17295 3455
rect 17255 3420 17260 3450
rect 17290 3420 17295 3450
rect 17255 3415 17295 3420
rect 17435 3450 17475 3455
rect 17435 3420 17440 3450
rect 17470 3420 17475 3450
rect 17435 3415 17475 3420
rect 17615 3450 17655 3455
rect 17615 3420 17620 3450
rect 17650 3420 17655 3450
rect 17615 3415 17655 3420
rect 17795 3450 17835 3455
rect 17795 3420 17800 3450
rect 17830 3420 17835 3450
rect 17795 3415 17835 3420
rect 17975 3450 18015 3455
rect 17975 3420 17980 3450
rect 18010 3420 18015 3450
rect 17975 3415 18015 3420
rect 18155 3450 18195 3455
rect 18155 3420 18160 3450
rect 18190 3420 18195 3450
rect 18155 3415 18195 3420
rect 18335 3450 18375 3455
rect 18335 3420 18340 3450
rect 18370 3420 18375 3450
rect 18335 3415 18375 3420
rect 18515 3450 18555 3455
rect 18515 3420 18520 3450
rect 18550 3420 18555 3450
rect 18515 3415 18555 3420
rect 18695 3450 18735 3455
rect 18695 3420 18700 3450
rect 18730 3420 18735 3450
rect 18695 3415 18735 3420
rect 18875 3450 18915 3455
rect 18875 3420 18880 3450
rect 18910 3420 18915 3450
rect 18875 3415 18915 3420
rect 19055 3450 19095 3455
rect 19055 3420 19060 3450
rect 19090 3420 19095 3450
rect 19055 3415 19095 3420
rect 19235 3450 19275 3455
rect 19235 3420 19240 3450
rect 19270 3420 19275 3450
rect 19235 3415 19275 3420
rect 19415 3450 19455 3455
rect 19415 3420 19420 3450
rect 19450 3420 19455 3450
rect 19415 3415 19455 3420
rect 19595 3450 19635 3455
rect 19595 3420 19600 3450
rect 19630 3420 19635 3450
rect 19595 3415 19635 3420
rect 19775 3450 19815 3455
rect 19775 3420 19780 3450
rect 19810 3420 19815 3450
rect 19775 3415 19815 3420
rect 19955 3450 19995 3455
rect 19955 3420 19960 3450
rect 19990 3420 19995 3450
rect 19955 3415 19995 3420
rect 20675 3450 20715 3455
rect 20675 3420 20680 3450
rect 20710 3420 20715 3450
rect 20675 3415 20715 3420
rect 20810 3450 20850 4375
rect 20810 3420 20815 3450
rect 20845 3420 20850 3450
rect 20810 3415 20850 3420
<< via1 >>
rect 9160 4365 9190 4370
rect 9160 4345 9165 4365
rect 9165 4345 9185 4365
rect 9185 4345 9190 4365
rect 9160 4340 9190 4345
rect 9880 4365 9910 4370
rect 9880 4345 9885 4365
rect 9885 4345 9905 4365
rect 9905 4345 9910 4365
rect 9880 4340 9910 4345
rect 10060 4365 10090 4370
rect 10060 4345 10065 4365
rect 10065 4345 10085 4365
rect 10085 4345 10090 4365
rect 10060 4340 10090 4345
rect 10240 4365 10270 4370
rect 10240 4345 10245 4365
rect 10245 4345 10265 4365
rect 10265 4345 10270 4365
rect 10240 4340 10270 4345
rect 10420 4365 10450 4370
rect 10420 4345 10425 4365
rect 10425 4345 10445 4365
rect 10445 4345 10450 4365
rect 10420 4340 10450 4345
rect 10600 4365 10630 4370
rect 10600 4345 10605 4365
rect 10605 4345 10625 4365
rect 10625 4345 10630 4365
rect 10600 4340 10630 4345
rect 10780 4365 10810 4370
rect 10780 4345 10785 4365
rect 10785 4345 10805 4365
rect 10805 4345 10810 4365
rect 10780 4340 10810 4345
rect 10960 4365 10990 4370
rect 10960 4345 10965 4365
rect 10965 4345 10985 4365
rect 10985 4345 10990 4365
rect 10960 4340 10990 4345
rect 11140 4365 11170 4370
rect 11140 4345 11145 4365
rect 11145 4345 11165 4365
rect 11165 4345 11170 4365
rect 11140 4340 11170 4345
rect 11320 4365 11350 4370
rect 11320 4345 11325 4365
rect 11325 4345 11345 4365
rect 11345 4345 11350 4365
rect 11320 4340 11350 4345
rect 11500 4365 11530 4370
rect 11500 4345 11505 4365
rect 11505 4345 11525 4365
rect 11525 4345 11530 4365
rect 11500 4340 11530 4345
rect 11680 4365 11710 4370
rect 11680 4345 11685 4365
rect 11685 4345 11705 4365
rect 11705 4345 11710 4365
rect 11680 4340 11710 4345
rect 11860 4365 11890 4370
rect 11860 4345 11865 4365
rect 11865 4345 11885 4365
rect 11885 4345 11890 4365
rect 11860 4340 11890 4345
rect 12040 4365 12070 4370
rect 12040 4345 12045 4365
rect 12045 4345 12065 4365
rect 12065 4345 12070 4365
rect 12040 4340 12070 4345
rect 12220 4365 12250 4370
rect 12220 4345 12225 4365
rect 12225 4345 12245 4365
rect 12245 4345 12250 4365
rect 12220 4340 12250 4345
rect 12400 4365 12430 4370
rect 12400 4345 12405 4365
rect 12405 4345 12425 4365
rect 12425 4345 12430 4365
rect 12400 4340 12430 4345
rect 12580 4365 12610 4370
rect 12580 4345 12585 4365
rect 12585 4345 12605 4365
rect 12605 4345 12610 4365
rect 12580 4340 12610 4345
rect 12760 4365 12790 4370
rect 12760 4345 12765 4365
rect 12765 4345 12785 4365
rect 12785 4345 12790 4365
rect 12760 4340 12790 4345
rect 12940 4365 12970 4370
rect 12940 4345 12945 4365
rect 12945 4345 12965 4365
rect 12965 4345 12970 4365
rect 12940 4340 12970 4345
rect 13120 4365 13150 4370
rect 13120 4345 13125 4365
rect 13125 4345 13145 4365
rect 13145 4345 13150 4365
rect 13120 4340 13150 4345
rect 13300 4365 13330 4370
rect 13300 4345 13305 4365
rect 13305 4345 13325 4365
rect 13325 4345 13330 4365
rect 13300 4340 13330 4345
rect 13480 4365 13510 4370
rect 13480 4345 13485 4365
rect 13485 4345 13505 4365
rect 13505 4345 13510 4365
rect 13480 4340 13510 4345
rect 13660 4365 13690 4370
rect 13660 4345 13665 4365
rect 13665 4345 13685 4365
rect 13685 4345 13690 4365
rect 13660 4340 13690 4345
rect 13840 4365 13870 4370
rect 13840 4345 13845 4365
rect 13845 4345 13865 4365
rect 13865 4345 13870 4365
rect 13840 4340 13870 4345
rect 14020 4365 14050 4370
rect 14020 4345 14025 4365
rect 14025 4345 14045 4365
rect 14045 4345 14050 4365
rect 14020 4340 14050 4345
rect 14200 4365 14230 4370
rect 14200 4345 14205 4365
rect 14205 4345 14225 4365
rect 14225 4345 14230 4365
rect 14200 4340 14230 4345
rect 14380 4365 14410 4370
rect 14380 4345 14385 4365
rect 14385 4345 14405 4365
rect 14405 4345 14410 4365
rect 14380 4340 14410 4345
rect 14560 4365 14590 4370
rect 14560 4345 14565 4365
rect 14565 4345 14585 4365
rect 14585 4345 14590 4365
rect 14560 4340 14590 4345
rect 14740 4365 14770 4370
rect 14740 4345 14745 4365
rect 14745 4345 14765 4365
rect 14765 4345 14770 4365
rect 14740 4340 14770 4345
rect 14920 4365 14950 4370
rect 14920 4345 14925 4365
rect 14925 4345 14945 4365
rect 14945 4345 14950 4365
rect 14920 4340 14950 4345
rect 15100 4365 15130 4370
rect 15100 4345 15105 4365
rect 15105 4345 15125 4365
rect 15125 4345 15130 4365
rect 15100 4340 15130 4345
rect 15280 4365 15310 4370
rect 15280 4345 15285 4365
rect 15285 4345 15305 4365
rect 15305 4345 15310 4365
rect 15280 4340 15310 4345
rect 15460 4365 15490 4370
rect 15460 4345 15465 4365
rect 15465 4345 15485 4365
rect 15485 4345 15490 4365
rect 15460 4340 15490 4345
rect 15640 4365 15670 4370
rect 15640 4345 15645 4365
rect 15645 4345 15665 4365
rect 15665 4345 15670 4365
rect 15640 4340 15670 4345
rect 15820 4365 15850 4370
rect 15820 4345 15825 4365
rect 15825 4345 15845 4365
rect 15845 4345 15850 4365
rect 15820 4340 15850 4345
rect 16000 4365 16030 4370
rect 16000 4345 16005 4365
rect 16005 4345 16025 4365
rect 16025 4345 16030 4365
rect 16000 4340 16030 4345
rect 16180 4365 16210 4370
rect 16180 4345 16185 4365
rect 16185 4345 16205 4365
rect 16205 4345 16210 4365
rect 16180 4340 16210 4345
rect 16360 4365 16390 4370
rect 16360 4345 16365 4365
rect 16365 4345 16385 4365
rect 16385 4345 16390 4365
rect 16360 4340 16390 4345
rect 16540 4365 16570 4370
rect 16540 4345 16545 4365
rect 16545 4345 16565 4365
rect 16565 4345 16570 4365
rect 16540 4340 16570 4345
rect 16720 4365 16750 4370
rect 16720 4345 16725 4365
rect 16725 4345 16745 4365
rect 16745 4345 16750 4365
rect 16720 4340 16750 4345
rect 16900 4365 16930 4370
rect 16900 4345 16905 4365
rect 16905 4345 16925 4365
rect 16925 4345 16930 4365
rect 16900 4340 16930 4345
rect 17080 4365 17110 4370
rect 17080 4345 17085 4365
rect 17085 4345 17105 4365
rect 17105 4345 17110 4365
rect 17080 4340 17110 4345
rect 17260 4365 17290 4370
rect 17260 4345 17265 4365
rect 17265 4345 17285 4365
rect 17285 4345 17290 4365
rect 17260 4340 17290 4345
rect 17440 4365 17470 4370
rect 17440 4345 17445 4365
rect 17445 4345 17465 4365
rect 17465 4345 17470 4365
rect 17440 4340 17470 4345
rect 17620 4365 17650 4370
rect 17620 4345 17625 4365
rect 17625 4345 17645 4365
rect 17645 4345 17650 4365
rect 17620 4340 17650 4345
rect 17800 4365 17830 4370
rect 17800 4345 17805 4365
rect 17805 4345 17825 4365
rect 17825 4345 17830 4365
rect 17800 4340 17830 4345
rect 17980 4365 18010 4370
rect 17980 4345 17985 4365
rect 17985 4345 18005 4365
rect 18005 4345 18010 4365
rect 17980 4340 18010 4345
rect 18160 4365 18190 4370
rect 18160 4345 18165 4365
rect 18165 4345 18185 4365
rect 18185 4345 18190 4365
rect 18160 4340 18190 4345
rect 18340 4365 18370 4370
rect 18340 4345 18345 4365
rect 18345 4345 18365 4365
rect 18365 4345 18370 4365
rect 18340 4340 18370 4345
rect 18520 4365 18550 4370
rect 18520 4345 18525 4365
rect 18525 4345 18545 4365
rect 18545 4345 18550 4365
rect 18520 4340 18550 4345
rect 18700 4365 18730 4370
rect 18700 4345 18705 4365
rect 18705 4345 18725 4365
rect 18725 4345 18730 4365
rect 18700 4340 18730 4345
rect 18880 4365 18910 4370
rect 18880 4345 18885 4365
rect 18885 4345 18905 4365
rect 18905 4345 18910 4365
rect 18880 4340 18910 4345
rect 19060 4365 19090 4370
rect 19060 4345 19065 4365
rect 19065 4345 19085 4365
rect 19085 4345 19090 4365
rect 19060 4340 19090 4345
rect 19240 4365 19270 4370
rect 19240 4345 19245 4365
rect 19245 4345 19265 4365
rect 19265 4345 19270 4365
rect 19240 4340 19270 4345
rect 19420 4365 19450 4370
rect 19420 4345 19425 4365
rect 19425 4345 19445 4365
rect 19445 4345 19450 4365
rect 19420 4340 19450 4345
rect 19600 4365 19630 4370
rect 19600 4345 19605 4365
rect 19605 4345 19625 4365
rect 19625 4345 19630 4365
rect 19600 4340 19630 4345
rect 19780 4365 19810 4370
rect 19780 4345 19785 4365
rect 19785 4345 19805 4365
rect 19805 4345 19810 4365
rect 19780 4340 19810 4345
rect 19960 4365 19990 4370
rect 19960 4345 19965 4365
rect 19965 4345 19985 4365
rect 19985 4345 19990 4365
rect 19960 4340 19990 4345
rect 20680 4365 20710 4370
rect 20680 4345 20685 4365
rect 20685 4345 20705 4365
rect 20705 4345 20710 4365
rect 20680 4340 20710 4345
rect 9025 3445 9055 3450
rect 9025 3425 9030 3445
rect 9030 3425 9050 3445
rect 9050 3425 9055 3445
rect 9025 3420 9055 3425
rect 9160 3445 9190 3450
rect 9160 3425 9165 3445
rect 9165 3425 9185 3445
rect 9185 3425 9190 3445
rect 9160 3420 9190 3425
rect 9880 3445 9910 3450
rect 9880 3425 9885 3445
rect 9885 3425 9905 3445
rect 9905 3425 9910 3445
rect 9880 3420 9910 3425
rect 10060 3445 10090 3450
rect 10060 3425 10065 3445
rect 10065 3425 10085 3445
rect 10085 3425 10090 3445
rect 10060 3420 10090 3425
rect 10240 3445 10270 3450
rect 10240 3425 10245 3445
rect 10245 3425 10265 3445
rect 10265 3425 10270 3445
rect 10240 3420 10270 3425
rect 10420 3445 10450 3450
rect 10420 3425 10425 3445
rect 10425 3425 10445 3445
rect 10445 3425 10450 3445
rect 10420 3420 10450 3425
rect 10600 3445 10630 3450
rect 10600 3425 10605 3445
rect 10605 3425 10625 3445
rect 10625 3425 10630 3445
rect 10600 3420 10630 3425
rect 10780 3445 10810 3450
rect 10780 3425 10785 3445
rect 10785 3425 10805 3445
rect 10805 3425 10810 3445
rect 10780 3420 10810 3425
rect 10960 3445 10990 3450
rect 10960 3425 10965 3445
rect 10965 3425 10985 3445
rect 10985 3425 10990 3445
rect 10960 3420 10990 3425
rect 11140 3445 11170 3450
rect 11140 3425 11145 3445
rect 11145 3425 11165 3445
rect 11165 3425 11170 3445
rect 11140 3420 11170 3425
rect 11320 3445 11350 3450
rect 11320 3425 11325 3445
rect 11325 3425 11345 3445
rect 11345 3425 11350 3445
rect 11320 3420 11350 3425
rect 11500 3445 11530 3450
rect 11500 3425 11505 3445
rect 11505 3425 11525 3445
rect 11525 3425 11530 3445
rect 11500 3420 11530 3425
rect 11680 3445 11710 3450
rect 11680 3425 11685 3445
rect 11685 3425 11705 3445
rect 11705 3425 11710 3445
rect 11680 3420 11710 3425
rect 11860 3445 11890 3450
rect 11860 3425 11865 3445
rect 11865 3425 11885 3445
rect 11885 3425 11890 3445
rect 11860 3420 11890 3425
rect 12040 3445 12070 3450
rect 12040 3425 12045 3445
rect 12045 3425 12065 3445
rect 12065 3425 12070 3445
rect 12040 3420 12070 3425
rect 12220 3445 12250 3450
rect 12220 3425 12225 3445
rect 12225 3425 12245 3445
rect 12245 3425 12250 3445
rect 12220 3420 12250 3425
rect 12400 3445 12430 3450
rect 12400 3425 12405 3445
rect 12405 3425 12425 3445
rect 12425 3425 12430 3445
rect 12400 3420 12430 3425
rect 12580 3445 12610 3450
rect 12580 3425 12585 3445
rect 12585 3425 12605 3445
rect 12605 3425 12610 3445
rect 12580 3420 12610 3425
rect 12760 3445 12790 3450
rect 12760 3425 12765 3445
rect 12765 3425 12785 3445
rect 12785 3425 12790 3445
rect 12760 3420 12790 3425
rect 12940 3445 12970 3450
rect 12940 3425 12945 3445
rect 12945 3425 12965 3445
rect 12965 3425 12970 3445
rect 12940 3420 12970 3425
rect 13120 3445 13150 3450
rect 13120 3425 13125 3445
rect 13125 3425 13145 3445
rect 13145 3425 13150 3445
rect 13120 3420 13150 3425
rect 13300 3445 13330 3450
rect 13300 3425 13305 3445
rect 13305 3425 13325 3445
rect 13325 3425 13330 3445
rect 13300 3420 13330 3425
rect 13480 3445 13510 3450
rect 13480 3425 13485 3445
rect 13485 3425 13505 3445
rect 13505 3425 13510 3445
rect 13480 3420 13510 3425
rect 13660 3445 13690 3450
rect 13660 3425 13665 3445
rect 13665 3425 13685 3445
rect 13685 3425 13690 3445
rect 13660 3420 13690 3425
rect 13840 3445 13870 3450
rect 13840 3425 13845 3445
rect 13845 3425 13865 3445
rect 13865 3425 13870 3445
rect 13840 3420 13870 3425
rect 14020 3445 14050 3450
rect 14020 3425 14025 3445
rect 14025 3425 14045 3445
rect 14045 3425 14050 3445
rect 14020 3420 14050 3425
rect 14200 3445 14230 3450
rect 14200 3425 14205 3445
rect 14205 3425 14225 3445
rect 14225 3425 14230 3445
rect 14200 3420 14230 3425
rect 14380 3445 14410 3450
rect 14380 3425 14385 3445
rect 14385 3425 14405 3445
rect 14405 3425 14410 3445
rect 14380 3420 14410 3425
rect 14560 3445 14590 3450
rect 14560 3425 14565 3445
rect 14565 3425 14585 3445
rect 14585 3425 14590 3445
rect 14560 3420 14590 3425
rect 14740 3445 14770 3450
rect 14740 3425 14745 3445
rect 14745 3425 14765 3445
rect 14765 3425 14770 3445
rect 14740 3420 14770 3425
rect 14920 3445 14950 3450
rect 14920 3425 14925 3445
rect 14925 3425 14945 3445
rect 14945 3425 14950 3445
rect 14920 3420 14950 3425
rect 15100 3445 15130 3450
rect 15100 3425 15105 3445
rect 15105 3425 15125 3445
rect 15125 3425 15130 3445
rect 15100 3420 15130 3425
rect 15280 3445 15310 3450
rect 15280 3425 15285 3445
rect 15285 3425 15305 3445
rect 15305 3425 15310 3445
rect 15280 3420 15310 3425
rect 15460 3445 15490 3450
rect 15460 3425 15465 3445
rect 15465 3425 15485 3445
rect 15485 3425 15490 3445
rect 15460 3420 15490 3425
rect 15640 3445 15670 3450
rect 15640 3425 15645 3445
rect 15645 3425 15665 3445
rect 15665 3425 15670 3445
rect 15640 3420 15670 3425
rect 15820 3445 15850 3450
rect 15820 3425 15825 3445
rect 15825 3425 15845 3445
rect 15845 3425 15850 3445
rect 15820 3420 15850 3425
rect 16000 3445 16030 3450
rect 16000 3425 16005 3445
rect 16005 3425 16025 3445
rect 16025 3425 16030 3445
rect 16000 3420 16030 3425
rect 16180 3445 16210 3450
rect 16180 3425 16185 3445
rect 16185 3425 16205 3445
rect 16205 3425 16210 3445
rect 16180 3420 16210 3425
rect 16360 3445 16390 3450
rect 16360 3425 16365 3445
rect 16365 3425 16385 3445
rect 16385 3425 16390 3445
rect 16360 3420 16390 3425
rect 16540 3445 16570 3450
rect 16540 3425 16545 3445
rect 16545 3425 16565 3445
rect 16565 3425 16570 3445
rect 16540 3420 16570 3425
rect 16720 3445 16750 3450
rect 16720 3425 16725 3445
rect 16725 3425 16745 3445
rect 16745 3425 16750 3445
rect 16720 3420 16750 3425
rect 16900 3445 16930 3450
rect 16900 3425 16905 3445
rect 16905 3425 16925 3445
rect 16925 3425 16930 3445
rect 16900 3420 16930 3425
rect 17080 3445 17110 3450
rect 17080 3425 17085 3445
rect 17085 3425 17105 3445
rect 17105 3425 17110 3445
rect 17080 3420 17110 3425
rect 17260 3445 17290 3450
rect 17260 3425 17265 3445
rect 17265 3425 17285 3445
rect 17285 3425 17290 3445
rect 17260 3420 17290 3425
rect 17440 3445 17470 3450
rect 17440 3425 17445 3445
rect 17445 3425 17465 3445
rect 17465 3425 17470 3445
rect 17440 3420 17470 3425
rect 17620 3445 17650 3450
rect 17620 3425 17625 3445
rect 17625 3425 17645 3445
rect 17645 3425 17650 3445
rect 17620 3420 17650 3425
rect 17800 3445 17830 3450
rect 17800 3425 17805 3445
rect 17805 3425 17825 3445
rect 17825 3425 17830 3445
rect 17800 3420 17830 3425
rect 17980 3445 18010 3450
rect 17980 3425 17985 3445
rect 17985 3425 18005 3445
rect 18005 3425 18010 3445
rect 17980 3420 18010 3425
rect 18160 3445 18190 3450
rect 18160 3425 18165 3445
rect 18165 3425 18185 3445
rect 18185 3425 18190 3445
rect 18160 3420 18190 3425
rect 18340 3445 18370 3450
rect 18340 3425 18345 3445
rect 18345 3425 18365 3445
rect 18365 3425 18370 3445
rect 18340 3420 18370 3425
rect 18520 3445 18550 3450
rect 18520 3425 18525 3445
rect 18525 3425 18545 3445
rect 18545 3425 18550 3445
rect 18520 3420 18550 3425
rect 18700 3445 18730 3450
rect 18700 3425 18705 3445
rect 18705 3425 18725 3445
rect 18725 3425 18730 3445
rect 18700 3420 18730 3425
rect 18880 3445 18910 3450
rect 18880 3425 18885 3445
rect 18885 3425 18905 3445
rect 18905 3425 18910 3445
rect 18880 3420 18910 3425
rect 19060 3445 19090 3450
rect 19060 3425 19065 3445
rect 19065 3425 19085 3445
rect 19085 3425 19090 3445
rect 19060 3420 19090 3425
rect 19240 3445 19270 3450
rect 19240 3425 19245 3445
rect 19245 3425 19265 3445
rect 19265 3425 19270 3445
rect 19240 3420 19270 3425
rect 19420 3445 19450 3450
rect 19420 3425 19425 3445
rect 19425 3425 19445 3445
rect 19445 3425 19450 3445
rect 19420 3420 19450 3425
rect 19600 3445 19630 3450
rect 19600 3425 19605 3445
rect 19605 3425 19625 3445
rect 19625 3425 19630 3445
rect 19600 3420 19630 3425
rect 19780 3445 19810 3450
rect 19780 3425 19785 3445
rect 19785 3425 19805 3445
rect 19805 3425 19810 3445
rect 19780 3420 19810 3425
rect 19960 3445 19990 3450
rect 19960 3425 19965 3445
rect 19965 3425 19985 3445
rect 19985 3425 19990 3445
rect 19960 3420 19990 3425
rect 20680 3445 20710 3450
rect 20680 3425 20685 3445
rect 20685 3425 20705 3445
rect 20705 3425 20710 3445
rect 20680 3420 20710 3425
rect 20815 3445 20845 3450
rect 20815 3425 20820 3445
rect 20820 3425 20840 3445
rect 20840 3425 20845 3445
rect 20815 3420 20845 3425
<< metal2 >>
rect 9155 4370 20720 4375
rect 9155 4340 9160 4370
rect 9190 4340 9880 4370
rect 9910 4340 10060 4370
rect 10090 4340 10240 4370
rect 10270 4340 10420 4370
rect 10450 4340 10600 4370
rect 10630 4340 10780 4370
rect 10810 4340 10960 4370
rect 10990 4340 11140 4370
rect 11170 4340 11320 4370
rect 11350 4340 11500 4370
rect 11530 4340 11680 4370
rect 11710 4340 11860 4370
rect 11890 4340 12040 4370
rect 12070 4340 12220 4370
rect 12250 4340 12400 4370
rect 12430 4340 12580 4370
rect 12610 4340 12760 4370
rect 12790 4340 12940 4370
rect 12970 4340 13120 4370
rect 13150 4340 13300 4370
rect 13330 4340 13480 4370
rect 13510 4340 13660 4370
rect 13690 4340 13840 4370
rect 13870 4340 14020 4370
rect 14050 4340 14200 4370
rect 14230 4340 14380 4370
rect 14410 4340 14560 4370
rect 14590 4340 14740 4370
rect 14770 4340 14920 4370
rect 14950 4340 15100 4370
rect 15130 4340 15280 4370
rect 15310 4340 15460 4370
rect 15490 4340 15640 4370
rect 15670 4340 15820 4370
rect 15850 4340 16000 4370
rect 16030 4340 16180 4370
rect 16210 4340 16360 4370
rect 16390 4340 16540 4370
rect 16570 4340 16720 4370
rect 16750 4340 16900 4370
rect 16930 4340 17080 4370
rect 17110 4340 17260 4370
rect 17290 4340 17440 4370
rect 17470 4340 17620 4370
rect 17650 4340 17800 4370
rect 17830 4340 17980 4370
rect 18010 4340 18160 4370
rect 18190 4340 18340 4370
rect 18370 4340 18520 4370
rect 18550 4340 18700 4370
rect 18730 4340 18880 4370
rect 18910 4340 19060 4370
rect 19090 4340 19240 4370
rect 19270 4340 19420 4370
rect 19450 4340 19600 4370
rect 19630 4340 19780 4370
rect 19810 4340 19960 4370
rect 19990 4340 20680 4370
rect 20710 4340 20720 4370
rect 9155 4335 20720 4340
rect 9020 3450 20850 3455
rect 9020 3420 9025 3450
rect 9055 3420 9160 3450
rect 9190 3420 9880 3450
rect 9910 3420 10060 3450
rect 10090 3420 10240 3450
rect 10270 3420 10420 3450
rect 10450 3420 10600 3450
rect 10630 3420 10780 3450
rect 10810 3420 10960 3450
rect 10990 3420 11140 3450
rect 11170 3420 11320 3450
rect 11350 3420 11500 3450
rect 11530 3420 11680 3450
rect 11710 3420 11860 3450
rect 11890 3420 12040 3450
rect 12070 3420 12220 3450
rect 12250 3420 12400 3450
rect 12430 3420 12580 3450
rect 12610 3420 12760 3450
rect 12790 3420 12940 3450
rect 12970 3420 13120 3450
rect 13150 3420 13300 3450
rect 13330 3420 13480 3450
rect 13510 3420 13660 3450
rect 13690 3420 13840 3450
rect 13870 3420 14020 3450
rect 14050 3420 14200 3450
rect 14230 3420 14380 3450
rect 14410 3420 14560 3450
rect 14590 3420 14740 3450
rect 14770 3420 14920 3450
rect 14950 3420 15100 3450
rect 15130 3420 15280 3450
rect 15310 3420 15460 3450
rect 15490 3420 15640 3450
rect 15670 3420 15820 3450
rect 15850 3420 16000 3450
rect 16030 3420 16180 3450
rect 16210 3420 16360 3450
rect 16390 3420 16540 3450
rect 16570 3420 16720 3450
rect 16750 3420 16900 3450
rect 16930 3420 17080 3450
rect 17110 3420 17260 3450
rect 17290 3420 17440 3450
rect 17470 3420 17620 3450
rect 17650 3420 17800 3450
rect 17830 3420 17980 3450
rect 18010 3420 18160 3450
rect 18190 3420 18340 3450
rect 18370 3420 18520 3450
rect 18550 3420 18700 3450
rect 18730 3420 18880 3450
rect 18910 3420 19060 3450
rect 19090 3420 19240 3450
rect 19270 3420 19420 3450
rect 19450 3420 19600 3450
rect 19630 3420 19780 3450
rect 19810 3420 19960 3450
rect 19990 3420 20680 3450
rect 20710 3420 20815 3450
rect 20845 3420 20850 3450
rect 9020 3415 20850 3420
<< labels >>
rlabel metal2 9160 3435 9160 3435 1 VSSA
port 2 n
rlabel metal2 9160 4355 9160 4355 1 VDDA
port 1 n
rlabel locali 9165 3855 9165 3855 1 in
port 7 n
rlabel locali 9165 3975 9165 3975 1 p2
port 4 n
rlabel locali 9165 4015 9165 4015 1 p1
port 3 n
rlabel locali 9165 3695 9165 3695 1 n1
port 6 n
rlabel locali 9165 3735 9165 3735 1 n2
port 5 n
rlabel locali 9165 3895 9165 3895 1 out
port 8 n
rlabel locali 9165 3775 9165 3775 1 p3
rlabel locali 9165 4095 9165 4095 1 n3
rlabel locali 9165 3935 9165 3935 1 xp
rlabel locali 9165 3815 9165 3815 1 xn
<< end >>
