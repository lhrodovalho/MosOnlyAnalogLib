* NGSPICE file created from opamp.ext - technology: sky130A

.subckt ota VDDA VSSA P1 P2 N2 N1 INP INM OUT
X0 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.4e+12p pd=3.36e+07u as=5.2e+12p ps=7.28e+07u w=1e+06u l=500000u
X1 a_n1395_50# N2 OUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=6e+11p ps=8.4e+06u w=1e+06u l=500000u
X2 a_n5805_50# a_n6485_35# a_n5895_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X3 a_n8055_1845# N1 a_n8145_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X4 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2.4e+12p pd=3.36e+07u as=0p ps=0u w=1e+06u l=500000u
X5 OUT a_n6485_35# a_n4455_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X6 a_n1575_830# P2 a_n1665_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X7 a_n9225_1065# Z a_n9315_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X8 a_n9585_50# a_n10085_35# a_n9675_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X9 VDDA P1 a_n7335_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.4e+12p pd=1.96e+07u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X10 a_n11525_1795# a_n11525_1795# a_n11385_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=2e+11p pd=2.8e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X11 a_n5895_1845# a_n7205_1795# a_n5985_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X12 a_n725_35# a_n725_35# a_n405_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=2e+11p pd=2.8e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X13 a_n1395_1065# P2 X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X14 a_n4995_1845# N2 OUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X15 a_n725_1050# a_n725_1050# a_n585_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2e+11p pd=2.8e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X16 a_n10215_830# P2 a_n10305_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X17 a_n11205_50# a_n11525_35# a_n11525_35# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=2e+11p ps=2.8e+06u w=1e+06u l=500000u
X18 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X19 a_n3195_1845# a_n3605_1795# a_n3285_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X20 VSSA N1 a_n855_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1.4e+12p pd=1.96e+07u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X21 a_n2115_830# Z VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X22 a_n9765_1065# P2 a_n9855_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X23 a_n1935_50# N1 a_n2025_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X24 VDDA a_n725_780# a_n135_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X25 VSSA N1 a_n855_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X26 a_n7785_830# P2 a_n7875_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X27 a_n5985_50# a_n6485_35# a_n6075_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X28 a_n6435_1845# a_n7205_1795# a_n6525_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X29 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X30 a_n5535_1845# a_n7205_1795# a_n5625_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X31 a_n10755_830# P1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X32 a_n1035_1065# P1 a_n1125_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X33 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X34 a_n4905_50# a_n6485_35# a_n4995_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X35 a_n4545_50# a_n6485_35# a_n4635_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X36 a_n3735_1845# N2 a_n3825_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X37 a_n8955_50# a_n10085_35# a_n10085_35# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X38 a_n2655_830# P2 a_n2745_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X39 a_n1305_1845# N2 a_n1395_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X40 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X41 a_n11475_1845# a_n11525_1795# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X42 a_n6075_1845# a_n7205_1795# a_n7205_1795# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X43 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X44 X P2 a_n7335_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X45 a_n1305_50# N2 a_n1395_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X46 a_n4275_1845# N1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X47 a_n9945_1845# N2 a_n10035_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X48 a_n7695_50# N2 a_n7785_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X49 OUT N2 a_n6615_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X50 a_n10215_1065# P2 a_n10305_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X51 YP N1 a_n9135_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=8e+11p pd=1.12e+07u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X52 a_n4545_1065# P1 a_n4635_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X53 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X54 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X55 a_n6615_1845# a_n7205_1795# a_n6705_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X56 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X57 VDDA a_n725_1050# a_n135_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X58 a_n7785_1065# P1 a_n7875_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X59 a_n4815_1845# N2 a_n4905_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X60 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X61 a_n10755_1065# Z VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X62 a_n9585_1845# N1 a_n9675_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X63 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X64 a_n725_1795# a_n725_1795# a_n405_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=2e+11p pd=2.8e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X65 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X66 OUT N2 a_n1575_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X67 a_n7155_1845# a_n7205_1795# OUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X68 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X69 a_n7065_50# N1 a_n7155_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X70 a_n8235_50# a_n10085_35# a_n8325_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X71 a_n675_830# a_n725_780# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X72 a_n8325_1065# P2 a_n8415_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X73 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X74 a_n10395_1845# N2 YM VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=8e+11p ps=1.12e+07u w=1e+06u l=500000u
X75 a_n4455_50# a_n6485_35# a_n4545_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X76 a_n4455_1845# N1 a_n4545_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X77 VDDA P1 a_n3735_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X78 a_n2295_1845# a_n3605_1795# a_n2385_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X79 a_n8865_1065# P2 a_n8955_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X80 a_n1215_830# P2 a_n1305_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X81 VDDA Z a_n8055_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X82 a_n6885_830# P1 a_n6975_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X83 a_n10935_1845# a_n11525_1795# a_n11025_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X84 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X85 a_n10035_1845# N2 OUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X86 a_n2025_50# N1 a_n2115_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X87 a_n3195_50# N2 YP VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X88 YP N2 a_n7695_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X89 a_n8775_50# a_n10085_35# a_n8865_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X90 a_n4185_830# P2 a_n4275_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X91 a_n9945_50# a_n10085_35# a_n10035_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X92 a_n2835_1845# a_n3605_1795# a_n2925_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X93 a_n1755_830# P2 a_n1845_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X94 VDDA Z a_n9495_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X95 a_n10035_50# a_n10085_35# Z VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=6e+11p ps=8.4e+06u w=1e+06u l=500000u
X96 a_n8505_1065# P2 a_n8595_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X97 a_n7425_830# P1 a_n7515_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X98 X P2 a_n6615_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X99 a_n10575_1845# N1 a_n10665_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X100 a_n5175_1845# a_n7205_1795# a_n5265_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X101 a_n675_1065# a_n725_1050# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X102 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X103 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X104 a_n3375_1845# a_n3605_1795# a_n3465_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X105 a_n5175_50# a_n6485_35# a_n5265_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X106 a_n6345_50# a_n6485_35# a_n6435_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X107 a_n2475_1845# a_n3605_1795# a_n3605_1795# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X108 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X109 a_n8145_1845# N1 a_n8235_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X110 YP N2 a_n2655_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X111 X P2 a_n3735_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X112 a_n3735_50# N1 a_n3825_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X113 a_n225_830# a_n725_780# a_n725_780# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=2e+11p ps=2.8e+06u w=1e+06u l=500000u
X114 a_n7065_830# P1 a_n7155_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X115 a_n11525_1795# a_n11525_1795# a_n11205_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X116 a_n9315_50# a_n10085_35# a_n9405_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X117 a_n5715_1845# a_n7205_1795# a_n5805_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X118 a_n1215_1065# P2 a_n1305_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X119 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X120 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X121 a_n3915_1845# N2 YP VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X122 a_n10575_50# N1 a_n10665_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X123 a_n3015_1845# a_n3605_1795# a_n3105_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X124 Z N2 a_n8775_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X125 a_n4185_1065# P1 a_n4275_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X126 a_n7605_830# P2 a_n7695_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X127 a_n6255_1845# a_n7205_1795# a_n6345_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X128 YM N1 a_n6975_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X129 a_n5715_50# a_n6485_35# a_n5805_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X130 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X131 a_n7425_1065# P2 a_n7515_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X132 a_n4275_50# N2 OUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X133 a_n3105_50# N2 a_n3195_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X134 VDDA a_n11525_780# a_n10935_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X135 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X136 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X137 a_n3555_1845# a_n3605_1795# Z VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X138 a_n9495_50# a_n10085_35# a_n9585_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X139 a_n9855_50# a_n10085_35# a_n9945_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X140 a_n9225_1845# N1 a_n9315_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X141 a_n225_50# a_n725_35# a_n725_35# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X142 a_n4725_1065# P2 a_n4815_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X143 a_n2745_830# P2 a_n2835_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X144 a_n9495_1065# Z a_n9585_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X145 a_n1395_1845# N2 Z VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X146 a_n11525_35# a_n11525_35# a_n11205_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X147 a_n725_1795# a_n725_1795# a_n585_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X148 a_n225_1065# a_n725_1050# a_n725_1050# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X149 a_n11385_830# a_n11525_780# a_n11475_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X150 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X151 a_n10485_830# P1 a_n10575_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X152 YM N1 a_n1935_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X153 a_n675_50# a_n725_35# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X154 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X155 YM N2 a_n9855_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X156 a_n6255_50# a_n6485_35# a_n6345_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X157 a_n7425_50# N1 a_n7515_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X158 a_n3285_830# Z a_n3375_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X159 a_n1935_1845# a_n3605_1795# a_n2025_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X160 a_n4815_50# a_n6485_35# a_n4905_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X161 a_n1035_1845# N1 YP VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X162 a_n855_830# Z a_n945_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X163 a_n7605_1065# P1 a_n7695_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X164 a_n11025_830# a_n11525_780# a_n11525_780# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=2e+11p ps=2.8e+06u w=1e+06u l=500000u
X165 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X166 VDDA a_n11525_1050# a_n10935_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X167 a_n3825_830# P1 a_n3915_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X168 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X169 a_n1575_1845# a_n3605_1795# a_n1665_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X170 a_n1215_50# N2 a_n1305_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X171 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X172 a_n2385_50# N1 a_n2475_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X173 OUT N2 a_n7335_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X174 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X175 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X176 a_n10215_1845# N2 a_n10305_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X177 a_n4545_1845# N1 a_n4635_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X178 a_n11385_1065# a_n11525_1050# a_n11475_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X179 a_n10395_50# N2 YP VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X180 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X181 a_n10485_1065# Z a_n10575_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X182 a_n3465_830# Z a_n3555_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X183 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X184 a_n2115_1845# a_n3605_1795# a_n2205_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X185 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X186 a_n7785_1845# N1 a_n7875_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X187 VSSA a_n725_1795# a_n135_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X188 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X189 a_n6705_830# P2 a_n6795_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X190 a_n10755_1845# N1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X191 a_n5355_1845# a_n7205_1795# a_n5445_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X192 a_n855_1065# P1 a_n945_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X193 a_n1755_50# N2 YM VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X194 Z N2 a_n3015_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X195 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X196 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X197 a_n11025_1065# a_n11525_1050# a_n11525_1050# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=2e+11p ps=2.8e+06u w=1e+06u l=500000u
X198 a_n6975_50# N1 a_n7065_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X199 a_n4005_830# P2 a_n4095_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X200 a_n8145_50# a_n10085_35# a_n8235_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X201 a_n2655_1845# a_n3605_1795# a_n2745_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X202 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X203 YP N2 a_n8415_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X204 a_n3825_1065# P2 a_n3915_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X205 a_n405_830# a_n725_780# a_n725_780# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X206 a_n1845_830# Z a_n1935_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X207 a_n10935_50# a_n11525_35# a_n11025_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X208 a_n8595_1065# P2 Z VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2e+11p ps=2.8e+06u w=1e+06u l=500000u
X209 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X210 a_n8865_1845# N2 a_n8955_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X211 VDDA P1 a_n4455_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X212 VSSA N1 a_n8055_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X213 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X214 a_n2385_830# Z a_n2475_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X215 a_n9135_1065# Z a_n9225_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X216 a_n7515_50# N1 YP VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X217 OUT P2 a_n1575_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=2e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X218 a_n8685_50# a_n10085_35# a_n8775_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X219 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X220 X P2 a_n10215_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X221 a_n10305_50# N2 a_n10395_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X222 VSSA N1 a_n9495_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X223 a_n4905_1065# P2 a_n4995_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X224 a_n8505_1845# N2 a_n8595_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X225 a_n4005_1065# P1 a_n4095_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X226 Z P2 a_n3015_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X227 a_n2025_830# Z a_n2115_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X228 a_n9675_1065# Z a_n9765_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X229 a_n675_1845# a_n725_1795# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X230 a_n7695_830# P2 a_n7785_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X231 a_n5085_50# a_n6485_35# a_n5175_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X232 a_n405_1065# a_n725_1050# a_n725_1050# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X233 a_n6345_1845# a_n7205_1795# a_n6435_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X234 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X235 a_n2475_50# N1 YP VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X236 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X237 a_n10665_830# P1 a_n10755_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X238 VSSA N1 a_n3735_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X239 Z N2 a_n3735_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X240 a_n8055_50# a_n10085_35# a_n8145_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X241 a_n9225_50# a_n10085_35# a_n9315_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X242 a_n2565_830# P2 a_n2655_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X243 a_n1215_1845# N2 a_n1305_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X244 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X245 YP N1 a_n10575_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X246 a_n6885_1845# a_n7205_1795# a_n6975_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X247 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X248 a_n5985_1845# a_n7205_1795# a_n6075_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X249 a_n11205_830# a_n11525_780# a_n11525_780# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X250 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X251 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X252 a_n4185_1845# N1 a_n4275_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X253 a_n5625_50# a_n6485_35# a_n5715_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X254 OUT P2 a_n10215_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X255 a_n6795_50# N2 YM VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X256 a_n3105_830# P2 a_n3195_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X257 a_n1755_1845# a_n3605_1795# a_n1845_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X258 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X259 a_n3015_50# N2 a_n3105_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X260 a_n7425_1845# N2 a_n7515_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X261 a_n4185_50# N2 a_n4275_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X262 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X263 a_n6525_1845# a_n7205_1795# a_n6615_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X264 a_n9765_50# a_n10085_35# a_n9855_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X265 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X266 a_n945_830# Z a_n1035_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X267 a_n135_50# a_n725_35# a_n225_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X268 a_n7695_1065# P1 a_n7785_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X269 YM N2 a_n4815_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X270 a_n11025_50# a_n11525_35# a_n11525_35# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X271 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X272 a_n10665_1065# Z a_n10755_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X273 a_n9495_1845# N1 a_n9585_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X274 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X275 a_n225_1845# a_n725_1795# a_n725_1795# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X276 a_n7065_1845# a_n7205_1795# a_n7155_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X277 a_n585_50# a_n725_35# a_n675_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X278 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X279 a_n6165_50# a_n6485_35# a_n6255_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X280 a_n7335_50# N1 a_n7425_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X281 a_n585_830# a_n725_780# a_n675_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X282 a_n8235_1065# Z a_n8325_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X283 a_n3555_50# N1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X284 a_n4725_50# a_n6485_35# a_n4815_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X285 a_n11205_1065# a_n11525_1050# a_n11525_1050# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X286 X INM YM VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X287 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X288 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X289 YM N1 a_n7695_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X290 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X291 a_n8775_1065# P2 a_n8865_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X292 a_n1125_830# P2 a_n1215_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X293 a_n6795_830# P2 a_n6885_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X294 VSSA a_n11525_1795# a_n10935_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X295 a_n5445_1845# a_n7205_1795# a_n5535_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X296 a_n945_1065# P1 a_n1035_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X297 YM N2 a_n1215_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X298 a_n2295_50# N1 a_n2385_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X299 a_n6705_50# N2 a_n6795_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X300 a_n7875_50# N2 Z VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X301 a_n4095_830# P2 a_n4185_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X302 a_n2745_1845# a_n3605_1795# a_n2835_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X303 a_n1665_830# P2 a_n1755_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X304 a_n9315_1065# Z VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X305 a_n7335_830# P1 a_n7425_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X306 a_n11385_1845# a_n11525_1795# a_n11475_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X307 YM N1 a_n10575_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X308 OUT a_n7205_1795# a_n5175_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X309 a_n585_1065# a_n725_1050# a_n675_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X310 a_n10305_830# P2 a_n10395_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X311 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X312 a_n3285_1845# a_n3605_1795# a_n3375_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X313 a_n6485_35# a_n6485_35# a_n5535_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X314 a_n1665_50# N2 a_n1755_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X315 VDDA Z a_n2295_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X316 a_n9855_1065# P2 a_n9945_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X317 a_n2835_50# N2 Z VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X318 a_n135_830# a_n725_780# a_n225_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X319 a_n8955_1065# P2 a_n9045_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X320 a_n855_1845# N1 a_n945_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X321 a_n7875_830# P2 X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X322 a_n6975_830# P1 a_n7065_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X323 a_n8415_50# a_n10085_35# a_n8505_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X324 a_n11025_1845# a_n11525_1795# a_n11525_1795# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X325 a_n5625_1845# a_n7205_1795# a_n5715_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X326 a_n1125_1065# P2 a_n1215_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X327 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X328 a_n3825_1845# N2 a_n3915_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X329 VSSA a_n11525_35# a_n10935_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X330 a_n8595_1845# N2 Z VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X331 a_n4095_1065# P1 a_n4185_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X332 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X333 a_n7515_830# P1 a_n7605_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X334 a_n7205_1795# a_n7205_1795# a_n6255_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X335 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X336 a_n7335_1065# P2 a_n7425_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X337 VSSA N1 a_n2295_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X338 VSSA N1 a_n4455_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X339 a_n3375_50# N1 a_n3465_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X340 a_n3465_1845# a_n3605_1795# a_n3555_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X341 a_n8595_50# a_n10085_35# a_n8685_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X342 a_n10305_1065# P2 a_n10395_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X343 a_n9135_1845# N1 a_n9225_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X344 a_n4635_1065# P1 a_n4725_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X345 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X346 a_n10215_50# N2 a_n10305_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X347 a_n6705_1845# a_n7205_1795# a_n6795_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X348 a_n11385_50# a_n11525_35# a_n11475_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X349 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X350 a_n135_1065# a_n725_1050# a_n225_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X351 a_n7875_1065# P1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X352 a_n11525_780# a_n11525_780# a_n11385_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X353 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X354 a_n4905_1845# N2 a_n4995_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X355 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X356 YP N1 a_n4095_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X357 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X358 a_n945_50# N1 a_n1035_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X359 a_n9675_1845# N1 YM VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X360 a_n5355_50# a_n6485_35# a_n6485_35# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X361 a_n4995_50# a_n6485_35# a_n5085_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X362 a_n405_1845# a_n725_1795# a_n725_1795# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X363 a_n3195_830# P2 a_n3285_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X364 a_n1845_1845# a_n3605_1795# a_n1935_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X365 a_n3915_50# N1 YM VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X366 Z a_n10085_35# a_n8055_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X367 a_n9135_50# a_n10085_35# a_n9225_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X368 VDDA Z a_n855_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X369 a_n8415_1065# P2 a_n8505_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X370 a_n7515_1065# P2 a_n7605_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X371 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X372 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X373 a_n10755_50# N1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X374 a_n3735_830# P1 a_n3825_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X375 a_n2385_1845# a_n3605_1795# a_n2475_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X376 Z a_n3605_1795# a_n1575_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X377 a_n1305_830# P2 a_n1395_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X378 a_n5535_50# a_n6485_35# a_n5625_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X379 a_n8055_1065# Z a_n8145_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X380 a_n11475_830# a_n11525_780# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X381 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X382 OUT N2 a_n10215_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X383 a_n4095_50# N2 a_n4185_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X384 a_n8505_50# a_n10085_35# a_n8595_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X385 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X386 a_n11525_1050# a_n11525_1050# a_n11385_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X387 a_n9675_50# a_n10085_35# a_n9765_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X388 a_n4275_830# P2 X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X389 a_n4995_1065# P2 X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X390 a_n2925_1845# a_n3605_1795# a_n3015_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X391 a_n405_50# a_n725_35# a_n725_35# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X392 VSSA a_n725_35# a_n135_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X393 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X394 a_n2025_1845# a_n3605_1795# a_n2115_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X395 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X396 a_n7695_1845# N1 a_n7785_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X397 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X398 a_n6615_830# P2 a_n6705_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X399 a_n10665_1845# N1 a_n10755_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X400 a_n5265_1845# a_n7205_1795# a_n5355_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X401 VDDA P1 a_n855_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X402 a_n855_50# N1 a_n945_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X403 a_n725_35# a_n725_35# a_n585_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X404 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X405 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X406 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X407 a_n6075_50# a_n6485_35# a_n6165_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X408 VSSA N1 a_n7335_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X409 a_n3605_1795# a_n3605_1795# a_n2655_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X410 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X411 a_n8235_1845# N1 YP VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X412 a_n3465_50# N1 a_n3555_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X413 a_n3735_1065# P2 a_n3825_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X414 a_n4635_50# a_n6485_35# a_n4725_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X415 a_n725_780# a_n725_780# a_n405_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X416 a_n7155_830# P1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X417 a_n11205_1845# a_n11525_1795# a_n11525_1795# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X418 a_n5805_1845# a_n7205_1795# a_n5895_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X419 a_n1305_1065# P2 a_n1395_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X420 a_n11475_1065# a_n11525_1050# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X421 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X422 a_n10395_830# P2 a_n10485_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X423 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X424 a_n11475_50# a_n11525_35# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X425 a_n3105_1845# a_n3605_1795# a_n3195_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X426 a_n8775_1845# N2 a_n8865_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X427 a_n4275_1065# P1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X428 a_n1035_50# N1 YM VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X429 a_n2295_830# Z a_n2385_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X430 a_n9945_1065# P2 a_n10035_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X431 a_n9045_1065# Z a_n9135_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X432 a_n945_1845# N1 a_n1035_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X433 a_n6615_50# N2 a_n6705_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X434 a_n7785_50# N2 a_n7875_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X435 YM N2 a_n4095_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X436 a_n10935_830# a_n11525_780# a_n11025_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X437 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X438 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X439 a_n9315_1845# N1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X440 a_n4815_1065# P2 a_n4905_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X441 a_n2835_830# P2 Z VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X442 a_n9585_1065# Z a_n9675_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X443 a_n585_1845# a_n725_1795# a_n675_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X444 a_n725_1050# a_n725_1050# a_n405_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X445 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X446 a_n1575_50# N2 a_n1665_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X447 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X448 a_n10575_830# P1 a_n10665_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X449 a_n2745_50# N2 a_n2835_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X450 a_n9855_1845# N2 a_n9945_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X451 a_n7155_50# N1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X452 a_n8955_1845# N2 YP VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X453 a_n8325_50# a_n10085_35# a_n8415_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X454 a_n10395_1065# P2 a_n10485_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X455 a_n3375_830# Z a_n3465_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X456 a_n4455_1065# P1 a_n4545_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X457 a_n2475_830# Z a_n2565_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X458 YP N2 a_n1215_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X459 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X460 a_n6795_1845# a_n7205_1795# a_n6885_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X461 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X462 a_n11525_780# a_n11525_780# a_n11205_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X463 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X464 a_n4095_1845# N1 a_n4185_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X465 a_n10935_1065# a_n11525_1050# a_n11025_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X466 a_n3915_830# P1 a_n4005_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X467 a_n10035_1065# P2 OUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X468 a_n5895_50# a_n6485_35# a_n5985_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X469 a_n3015_830# P2 a_n3105_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X470 a_n1665_1845# a_n3605_1795# a_n1755_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X471 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X472 a_n2115_50# N1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X473 a_n7335_1845# N2 a_n7425_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X474 YP N1 a_n3375_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X475 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X476 a_n8865_50# a_n10085_35# a_n8955_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X477 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X478 a_n10305_1845# N2 a_n10395_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X479 a_n4635_1845# N1 YM VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X480 Z N2 a_n10215_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X481 a_n11525_35# a_n11525_35# a_n11385_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X482 a_n10575_1065# Z a_n10665_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X483 a_n3555_830# Z VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X484 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X485 a_n2205_1845# a_n3605_1795# a_n2295_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X486 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X487 a_n7875_1845# N1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X488 a_n135_1845# a_n725_1795# a_n225_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X489 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X490 a_n6975_1845# a_n7205_1795# a_n7065_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X491 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X492 a_n5265_50# a_n6485_35# a_n5355_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X493 a_n1395_830# P2 OUT VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X494 a_n6435_50# a_n6485_35# OUT VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X495 a_n725_780# a_n725_780# a_n585_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X496 a_n8145_1065# Z a_n8235_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X497 a_n2655_50# N2 a_n2745_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X498 a_n3825_50# N1 a_n3915_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X499 a_n11525_1050# a_n11525_1050# a_n11205_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X500 YM INM X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X501 a_n9405_50# a_n10085_35# a_n9495_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X502 a_n10085_35# a_n10085_35# a_n9135_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X503 X INP YP VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X504 a_n8415_1845# N2 a_n8505_1845# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X505 a_n3915_1065# P2 a_n4005_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X506 a_n7515_1845# N2 YM VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X507 a_n1935_830# Z a_n2025_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X508 YP INP X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X509 a_n10665_50# N1 a_n10755_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X510 Z P2 a_n8775_1065# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X511 a_n1035_830# Z a_n1125_830# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
.ends

.subckt buffer VDDA VSSA p1 p2 n2 n1 in out m1_18540_6950# m1_18720_6950# a_18100_8090#
+ m1_18900_6950# xp
X0 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=8e+12p pd=5.6e+07u as=1.44e+13p ps=1.008e+08u w=2e+06u l=1e+06u
X1 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X2 a_30950_6950# n2 a_30770_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X3 a_30410_6950# n2 a_30230_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X4 xn n3 a_27170_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X5 a_26810_6950# n3 xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X6 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X7 a_25730_6950# n3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=6.8e+12p ps=4.76e+07u w=2e+06u l=1e+06u
X8 a_19610_6950# a_18430_6920# a_19430_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X9 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10 VSSA n3 a_22490_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X11 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12 a_38690_8430# p3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=6.8e+12p ps=4.76e+07u w=2e+06u l=1e+06u
X13 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.44e+13p pd=1.008e+08u as=8e+12p ps=5.6e+07u w=2e+06u l=1e+06u
X14 a_39770_8430# p3 xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X15 p3 in xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1.6e+12p pd=1.12e+07u as=0p ps=0u w=2e+06u l=1e+06u
X16 xp in p3 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X17 a_30050_8430# p3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X18 n3 p2 a_31850_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=8e+11p pd=5.6e+06u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X19 a_32570_8430# p1 a_32390_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X20 a_24290_8430# p3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X21 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X22 a_27890_8430# p2 n3 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X23 VDDA p1 a_28250_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X24 a_31490_8430# p1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X25 a_39770_6950# n3 xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X26 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X27 a_38690_6950# n3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X28 a_32570_6950# n3 xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X29 a_30050_6950# n1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X30 a_29510_6950# n2 a_29330_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X31 xn in n3 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.6e+12p ps=1.12e+07u w=2e+06u l=1e+06u
X32 a_31490_6950# n3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X33 a_28970_6950# n2 a_28790_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X34 VSSA n3 a_28250_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X35 n3 in xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X36 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X37 a_24290_6950# n3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X38 a_31850_8430# p2 a_31670_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X39 a_35450_8430# p3 xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X40 VDDA p3 a_23930_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X41 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X42 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X43 a_27170_8430# p1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X44 n3 p2 a_27530_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X45 a_28250_8430# p1 a_28070_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X46 xp p3 a_30050_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X47 p3 in xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X48 VDDA p3 a_31130_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X49 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X50 a_21050_8430# p3 xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X51 a_35450_6950# n3 xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X52 VSSA n3 a_23930_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X53 n3 in xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X54 VSSA n1 a_31130_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X55 a_30770_6950# n2 p3 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=8e+11p ps=5.6e+06u w=2e+06u l=1e+06u
X56 a_30230_6950# n1 a_30050_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X57 a_28250_6950# n3 xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X58 xn in n3 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X59 a_27170_6950# n3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X60 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X61 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X62 a_21050_6950# n3 xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X63 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X64 p3 in xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X65 VDDA p3 a_29690_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X66 a_32390_8430# p2 a_32210_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X67 a_32930_8430# p3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X68 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X69 a_34010_8430# p3 xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X70 xp p3 a_34370_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X71 xp p3 a_35810_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X72 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X73 VDDA p3 a_36890_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X74 xp p3 a_28610_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X75 a_18530_8430# a_18430_8330# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X76 a_19070_8430# a_18430_8330# a_18430_8330# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=8e+11p ps=5.6e+06u w=2e+06u l=1e+06u
X77 xp p3 a_21410_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X78 VSSA n3 a_36890_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X79 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X80 xn n3 a_35810_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X81 xn n3 a_34370_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X82 a_34010_6950# n3 xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X83 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X84 a_32930_6950# n3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X85 xn in n3 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X86 VSSA n1 a_29690_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X87 a_29330_6950# n2 p3 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X88 a_28790_6950# n1 a_28610_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X89 a_19070_6950# a_18430_6920# a_18430_6920# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=8e+11p ps=5.6e+06u w=2e+06u l=1e+06u
X90 a_18530_6950# a_18430_6920# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X91 xn n3 a_21410_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X92 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X93 a_32210_8430# p2 n3 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X94 VDDA p1 a_32570_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X95 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X96 a_35810_8430# p3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X97 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X98 a_28610_8430# p3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X99 xp in p3 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X100 a_31130_8430# p3 xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X101 a_31670_8430# p1 a_31490_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X102 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X103 a_21410_8430# p3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X104 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X105 VDDA p3 a_25370_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X106 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X107 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X108 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X109 a_35810_6950# n3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X110 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X111 VSSA n3 a_32570_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X112 n3 in xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X113 xn n3 a_31490_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X114 a_31130_6950# n1 a_30950_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X115 p3 n2 a_28970_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X116 a_28610_6950# n1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X117 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X118 VSSA n3 a_25370_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X119 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X120 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X121 a_21410_6950# n3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X122 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X123 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X124 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X125 a_34370_8430# p3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X126 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X127 a_36890_8430# p3 xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X128 xp p3 a_37250_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X129 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X130 VDDA p3 a_38330_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X131 a_40030_8330# a_40030_8330# a_40310_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=8e+11p pd=5.6e+06u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X132 a_41030_8430# a_40030_8330# a_40030_8330# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X133 a_29690_8430# p3 xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X134 a_18430_8330# a_18430_8330# a_18710_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X135 a_19430_8430# a_18430_8330# a_18430_8330# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X136 a_19970_8430# p3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X137 a_22490_8430# p3 xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X138 xp p3 a_22850_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X139 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X140 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X141 xp p3 a_19970_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X142 a_41030_6950# a_40030_6920# a_40030_6920# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=8e+11p ps=5.6e+06u w=2e+06u l=1e+06u
X143 a_40030_6920# a_40030_6920# a_40310_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X144 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X145 VSSA n3 a_38330_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X146 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X147 xn n3 a_37250_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X148 a_36890_6950# n3 xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X149 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X150 a_34370_6950# n3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X151 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X152 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X153 a_29690_6950# n1 a_29510_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X154 a_19430_6950# a_18430_6920# a_18430_6920# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X155 a_19970_6950# n3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=2e+06u l=1e+06u
X156 a_22490_6950# n3 xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X157 xn n3 a_22850_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X158 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X159 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X160 a_18430_6920# a_18430_6920# a_18710_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X161 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X162 xn n3 a_19970_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X163 xp p3 a_32930_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X164 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X165 VDDA p3 a_35450_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X166 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X167 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X168 a_37250_8430# p3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X169 a_40310_8430# a_40030_8330# a_40130_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X170 a_40030_8330# a_40030_8330# a_40670_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X171 a_18710_8430# a_18430_8330# a_18530_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X172 a_18430_8330# a_18430_8330# a_19070_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X173 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X174 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X175 a_22850_8430# p3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X176 a_25370_8430# p3 xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X177 xp p3 a_25730_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X178 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X179 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X180 VDDA p3 a_21050_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X181 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X182 a_40030_6920# a_40030_6920# a_40670_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X183 a_40310_6950# a_40030_6920# a_40130_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X184 a_37250_6950# n3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X185 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X186 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X187 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X188 VSSA n3 a_35450_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X189 xn n3 a_32930_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X190 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X191 a_22850_6950# n3 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X192 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X193 xn n3 a_25730_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X194 a_25370_6950# n3 xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X195 a_18710_6950# a_18430_6920# a_18530_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X196 a_18430_6920# a_18430_6920# a_19070_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X197 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X198 VSSA n3 a_21050_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X199 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X200 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X201 VDDA p3 a_39770_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X202 VDDA p3 a_34010_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X203 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X204 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X205 a_38330_8430# p3 xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X206 xp p3 a_38690_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X207 VDDA a_40030_8330# a_41210_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X208 a_28070_8430# p2 a_27890_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X209 VDDA a_18430_8330# a_19610_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X210 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X211 a_23930_8430# p3 xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X212 xp p3 a_24290_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X213 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X214 VDDA p3 a_26810_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X215 a_27530_8430# p2 a_27350_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X216 xp in p3 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X217 VSSA a_40030_6920# a_41210_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=2e+06u l=1e+06u
X218 VSSA n3 a_39770_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X219 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X220 xn n3 a_38690_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X221 a_38330_6950# n3 xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X222 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X223 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X224 VSSA n3 a_34010_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X225 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X226 a_23930_6950# n3 xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X227 p3 n2 a_30410_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X228 xn in n3 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X229 n3 in xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X230 VSSA n3 a_26810_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X231 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X232 xn n3 a_24290_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X233 VSSA a_18430_6920# a_19610_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X234 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X235 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X236 a_40130_8430# a_40030_8330# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X237 a_40670_8430# a_40030_8330# a_40030_8330# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X238 a_41210_8430# a_40030_8330# a_41030_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X239 xp in p3 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X240 a_19610_8430# a_18430_8330# a_19430_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X241 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X242 VDDA p3 a_22490_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X243 out out xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X244 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X245 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X246 a_25730_8430# p3 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X247 xp out out VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X248 a_26810_8430# p3 xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X249 a_27350_8430# p1 a_27170_8430# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X250 p3 in xp VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X251 a_41210_6950# a_40030_6920# a_41030_6950# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X252 a_40670_6950# a_40030_6920# a_40030_6920# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X253 a_40130_6950# a_40030_6920# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X254 xn out out VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X255 out out xn VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
.ends

.subckt bias VDDA VSSA P1 P2 N2 N1
X0 a_1900_50# X VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=2.4e+12p ps=3.36e+07u w=1e+06u l=500000u
X1 a_9280_990# P2 a_9190_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X2 Y Y a_8200_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=2e+11p pd=2.8e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X3 X P2 a_1360_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=5.6e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X4 a_550_750# P1 a_460_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X5 a_n310_700# a_n310_700# a_n170_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X6 N1 N1 a_6760_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=5.6e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X7 a_5860_1690# Y a_5770_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X8 a_9460_750# P2 a_9370_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X9 a_4240_990# P0 a_4150_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X10 a_8560_750# P2 P2 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=2e+11p ps=2.8e+06u w=1e+06u l=500000u
X11 a_1810_990# P2 a_1720_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X12 a_820_1690# N2 a_730_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X13 a_4420_750# P2 a_4330_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X14 a_8830_1690# X a_8740_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X15 a_6760_50# N1 a_6670_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X16 a_9820_990# P1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=2.6e+12p ps=3.64e+07u w=1e+06u l=500000u
X17 a_7930_50# N1 a_7840_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X18 a_6400_1690# N1 a_6310_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X19 a_10000_750# P1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X20 P1 N1 a_3700_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=5.6e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X21 a_4780_990# P0 a_4690_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X22 a_9100_750# P2 a_9010_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X23 a_2080_50# X a_1990_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X24 a_1360_1690# N2 a_1270_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X25 a_4960_750# P0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X26 P2 P2 a_2260_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X27 a_6940_750# P2 a_6850_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X28 a_4060_750# N1 N1 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X29 Z X a_9280_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=8e+11p pd=1.12e+07u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X30 a_4330_1690# N1 a_4240_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X31 a_7300_50# N1 a_7210_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X32 a_8470_50# N1 a_8380_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X33 a_370_990# P1 a_280_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X34 a_1900_1690# N1 a_1810_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X35 a_4600_750# P1 a_4510_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X36 a_10270_990# P2 a_10180_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X37 a_9910_1690# X a_9820_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X38 a_7480_750# P0 a_7390_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X39 a_6580_750# P0 a_6490_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X40 a_2620_50# Y Y VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X41 a_10450_750# P2 a_10360_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X42 a_3790_50# N1 a_3700_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X43 a_4870_1690# Y a_4780_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X44 a_2440_750# P2 a_2350_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X45 a_7840_990# P1 a_7750_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X46 a_6040_50# Y a_5950_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X47 a_10810_990# a_10670_975# a_10720_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X48 a_5410_990# P2 a_5320_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X49 a_8020_750# P2 a_7930_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X50 a_9550_1690# X a_9460_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X51 a_7120_750# P2 P1 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=2e+11p ps=2.8e+06u w=1e+06u l=500000u
X52 a_9010_50# N1 a_8920_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X53 a_2980_750# P1 a_2890_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X54 a_2080_750# P1 a_1990_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X55 a_7390_1690# N1 a_7300_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X56 a_8380_990# P2 Y VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=2e+11p ps=2.8e+06u w=1e+06u l=500000u
X57 a_460_1690# N2 a_370_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X58 a_10270_50# N2 a_10180_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X59 a_10360_1690# X a_10270_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X60 a_3160_50# X a_3070_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X61 VDDA P0 a_5860_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X62 a_4330_50# N1 a_4240_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X63 a_5050_990# P2 a_4960_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X64 a_3340_990# P0 a_3250_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X65 a_7660_750# P0 a_7570_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X66 VSSA a_n310_35# a_100_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X67 a_3520_750# P1 a_3430_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X68 VDDA P1 a_820_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X69 a_5410_50# Y a_5320_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X70 a_2620_750# P2 Y VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X71 a_8920_990# P1 a_8830_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X72 Z X a_7840_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X73 a_100_1690# a_n310_1640# a_10_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X74 a_10670_1640# a_10670_1640# a_10810_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X75 a_5500_1690# Y a_5410_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X76 VSSA N1 a_9100_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X77 a_3880_990# P2 P1 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X78 a_2890_1690# N1 a_2800_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X79 a_8200_750# P2 a_8110_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X80 Z X a_640_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X81 a_10810_50# a_10670_35# a_10720_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X82 a_1450_990# P2 a_1360_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X83 a_3160_750# P1 a_3070_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X84 N2 P2 a_460_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=4e+11p pd=5.6e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X85 a_8470_1690# Y a_8380_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X86 a_3700_50# N1 a_3610_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X87 a_6040_750# P0 a_5950_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X88 a_9460_990# P2 X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X89 a_n310_975# a_n310_975# a_n170_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X90 VSSA N1 a_4780_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X91 a_5140_750# P0 a_5050_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X92 a_8560_990# P2 a_8470_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X93 VSSA N1 a_7480_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X94 a_n260_750# a_n310_700# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X95 a_3430_1690# N1 a_3340_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X96 a_4420_990# P0 a_4330_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X97 a_5950_50# Y a_5860_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X98 P0 Y a_5500_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=2e+11p pd=2.8e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X99 a_1000_1690# N2 N2 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=2e+11p ps=2.8e+06u w=1e+06u l=500000u
X100 a_n310_35# a_n310_35# a_n170_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X101 a_3700_750# P2 a_3610_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X102 a_10000_990# P2 a_9910_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X103 VSSA X a_8920_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X104 a_8560_50# N1 a_8470_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X105 a_11080_750# a_10670_700# a_10990_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X106 a_8110_1690# Y a_8020_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X107 a_9730_50# N2 a_9640_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X108 a_5680_750# P2 P0 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=2e+11p ps=2.8e+06u w=1e+06u l=500000u
X109 a_9100_990# P1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X110 a_1270_50# X a_1180_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X111 a_2440_50# Y a_2350_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X112 a_3970_1690# N1 a_3880_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X113 a_1540_750# P2 X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X114 a_4960_990# P2 a_4870_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X115 VSSA N1 a_2980_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X116 a_640_750# P2 a_550_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X117 a_4060_990# P2 a_3970_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X118 a_6940_990# P2 N1 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X119 a_n170_1690# a_n310_1640# a_n260_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X120 a_100_50# a_n310_35# a_10_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X121 Z Y a_8560_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X122 a_6220_750# P0 a_6130_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X123 a_6130_50# Y a_6040_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X124 VSSA N1 a_4420_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X125 a_3610_1690# N1 a_3520_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X126 a_1180_750# P1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X127 a_7480_990# P1 a_7390_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X128 a_4600_990# P0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X129 a_6490_1690# N1 a_6400_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X130 a_9100_50# N1 a_9010_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X131 a_5590_1690# Y a_5500_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X132 VDDA P2 a_9100_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X133 a_6580_990# P2 a_6490_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X134 a_2980_50# X Z VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X135 VSSA X a_1720_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X136 VDDA P1 a_10360_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X137 a_2440_990# P2 P2 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X138 a_6760_750# P2 a_6670_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X139 a_1720_750# P1 a_1630_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X140 a_4150_1690# N1 a_4060_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X141 a_7030_1690# N1 a_6940_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X142 a_8020_990# P2 a_7930_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X143 a_7120_990# P2 a_7030_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X144 VSSA N1 a_6040_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X145 a_9730_750# P2 a_9640_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X146 a_6670_50# N1 a_6580_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X147 a_7840_50# N1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X148 P2 N1 a_1900_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=5.6e+06u as=0p ps=0u w=1e+06u l=500000u
X149 a_2980_990# P2 a_2890_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X150 a_7300_750# P2 a_7210_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X151 a_2080_990# P2 a_1990_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X152 a_1090_1690# N2 a_1000_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X153 a_4690_750# P1 a_4600_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X154 a_2350_50# Y a_2260_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X155 a_3520_50# N1 a_3430_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X156 a_10540_750# P1 a_10450_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X157 a_2260_750# P2 a_2170_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X158 N1 N1 a_6580_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=4e+11p pd=5.6e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X159 a_7660_990# P1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X160 a_2530_1690# N1 a_2440_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X161 a_3520_990# P2 a_3430_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X162 VSSA N2 a_1540_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X163 a_2620_990# P2 a_2530_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X164 a_9640_1690# X a_9550_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X165 a_7210_50# N1 a_7120_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X166 a_2800_750# P2 a_2710_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X167 a_280_750# LO VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X168 a_8380_50# N1 a_8290_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X169 a_10_1690# a_n310_1640# a_n310_1640# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X170 a_10180_750# P2 a_10090_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X171 a_7210_1690# N1 a_7120_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X172 a_8200_990# P2 a_8110_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X173 a_2170_1690# N1 a_2080_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X174 a_6040_990# P1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X175 a_3160_990# P0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X176 a_5140_990# P2 a_5050_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X177 a_n260_990# a_n310_975# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X178 a_10720_750# a_10670_700# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X179 a_5320_750# P2 a_5230_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X180 a_7750_1690# X a_7660_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X181 a_10_50# a_n310_35# a_n310_35# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X182 VSSA a_n310_1640# a_100_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X183 VSSA N1 a_7660_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X184 a_3700_990# P2 a_3610_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X185 P2 N1 a_2620_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X186 a_10990_1690# a_10670_1640# a_10670_1640# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X187 a_8920_50# N1 P2 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X188 Z X a_10000_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X189 a_11080_990# a_10670_975# a_10990_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X190 a_5680_990# P0 a_5590_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X191 a_8290_750# P2 a_8200_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X192 a_10180_50# N2 a_10090_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X193 a_1540_990# P1 a_1450_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X194 a_5860_750# P2 a_5770_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X195 a_640_990# P2 N2 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X196 a_3070_50# X a_2980_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X197 a_4240_50# N1 N1 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X198 a_3250_1690# N1 a_3160_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X199 a_460_50# X VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X200 a_820_750# P2 X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X201 P0 Y a_5140_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X202 VSSA N1 LO VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2e+11p ps=2.8e+06u w=1e+06u l=500000u
X203 a_5320_50# Y a_5230_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X204 a_8830_750# P2 a_8740_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X205 a_6220_990# P1 a_6130_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X206 a_6490_50# N1 a_6400_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X207 a_6400_750# P0 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X208 a_3790_750# P2 a_3700_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X209 a_1180_990# P2 a_1090_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X210 a_9460_50# N2 a_9370_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X211 a_9190_990# P1 a_9100_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X212 a_1000_50# X a_910_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X213 a_640_50# X a_550_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X214 a_1360_750# P2 a_1270_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X215 VSSA a_10670_1640# a_11080_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X216 a_6760_990# N1 N1 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X217 a_5770_1690# Y a_5680_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X218 a_10720_50# a_10670_35# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X219 a_9370_750# P1 a_9280_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X220 a_3610_50# N1 a_3520_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X221 a_4780_50# N1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X222 a_730_1690# N2 a_640_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X223 a_4330_750# P2 a_4240_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X224 a_1720_990# P2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X225 a_8740_1690# X Z VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X226 a_5860_50# Y a_5770_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X227 VDDA P1 a_9640_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X228 P1 N1 a_6940_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X229 a_1900_750# P1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X230 VDDA P1 a_9820_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X231 a_7300_990# P1 a_7210_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X232 a_6310_1690# N1 a_6220_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X233 a_4690_990# P0 a_4600_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X234 a_9640_50# N2 a_9550_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X235 a_10000_50# N2 N2 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X236 a_1180_50# X X VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2e+11p ps=2.8e+06u w=1e+06u l=500000u
X237 VDDA P1 a_4780_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X238 a_10540_990# LO VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X239 a_2260_990# P2 a_2170_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X240 a_1270_1690# N2 a_1180_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X241 a_9280_1690# X a_9190_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X242 N1 LO P1 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X243 N1 LO P1 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X244 a_4240_1690# N1 a_4150_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X245 N2 P2 a_9460_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X246 a_6400_50# N1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X247 a_280_990# P1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X248 a_1810_1690# N1 a_1720_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X249 a_2800_990# P2 a_2710_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X250 a_10180_990# P2 X VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X251 a_9820_1690# X X VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X252 a_7390_750# P2 a_7300_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X253 a_460_750# P1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X254 a_550_50# X a_460_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X255 Z Y a_2800_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X256 a_1720_50# X a_1630_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X257 a_10360_750# P2 N2 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X258 a_4780_1690# Y a_4690_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X259 a_2350_1690# N1 a_2260_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X260 a_10720_990# a_10670_975# VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X261 a_5320_990# P2 P0 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X262 a_7930_750# P2 a_7840_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X263 a_6580_50# N1 a_6490_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X264 a_10670_700# a_10670_700# a_10810_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X265 a_100_750# a_n310_700# a_10_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X266 a_5500_750# P2 a_5410_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X267 a_2890_750# P2 a_2800_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X268 Y P2 a_8200_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X269 a_370_1690# N2 a_280_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X270 a_9550_50# N2 a_9460_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X271 a_10540_50# N2 a_10450_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X272 a_10270_1690# X a_10180_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X273 a_2260_50# Y Z VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X274 P2 P2 a_8380_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X275 a_5860_990# P0 a_5770_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X276 a_3430_50# N1 a_3340_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X277 a_7570_750# P0 a_7480_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X278 a_3430_750# P1 a_3340_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X279 a_820_990# P1 a_730_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X280 a_8830_990# P1 a_8740_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X281 a_7840_1690# X a_7750_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X282 a_1000_750# P1 a_910_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X283 a_10810_1690# a_10670_1640# a_10720_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X284 a_5410_1690# Y a_5320_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X285 a_7120_50# N1 P1 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X286 a_9010_750# P2 a_8920_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X287 a_6400_990# P2 a_6310_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X288 P1 P2 a_3700_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X289 a_8290_50# N1 a_8200_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X290 a_8110_750# P2 a_8020_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X291 N1 P2 a_3880_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X292 a_1360_990# P2 N2 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X293 a_3070_750# P1 a_2980_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X294 a_8380_1690# Y Y VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X295 a_2800_50# Y a_2710_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X296 X P2 a_9280_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X297 N1 N1 a_3880_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X298 a_n170_750# a_n310_700# a_n260_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X299 a_3340_1690# N1 a_3250_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X300 VSSA Y a_5860_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X301 a_4330_990# P0 a_4240_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X302 a_5050_1690# Y a_4960_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X303 a_8650_750# P2 a_8560_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X304 a_1900_990# P2 a_1810_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X305 N2 N2 a_820_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X306 a_4510_750# P2 a_4420_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X307 a_3610_750# P1 a_3520_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X308 a_8920_1690# X a_8830_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X309 a_7660_50# N1 a_7570_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X310 a_6490_750# P0 a_6400_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X311 a_9910_990# P1 a_9820_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X312 P2 N1 a_8740_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X313 P0 P2 a_5500_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X314 a_1540_50# X Z VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X315 a_3880_1690# N1 P1 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X316 a_4870_990# P0 a_4780_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X317 a_10090_50# N2 a_10000_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X318 a_10450_50# N2 a_10360_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X319 a_4510_50# N1 a_4420_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X320 a_1450_1690# N2 a_1360_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X321 a_n310_1640# a_n310_1640# a_n170_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X322 a_550_1690# N2 a_460_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X323 P1 P2 a_6940_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X324 N1 N1 a_4060_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X325 a_9460_1690# X Z VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X326 VSSA N1 LO VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X327 a_8560_1690# Y a_8470_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X328 a_6130_750# P0 a_6040_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X329 a_9550_990# P2 a_9460_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X330 a_5230_50# Y a_5140_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X331 a_1990_750# P1 a_1900_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X332 a_4420_1690# N1 a_4330_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X333 VDDA P1 a_1000_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X334 a_7390_990# P1 a_7300_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X335 a_8200_50# N1 P2 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X336 a_9370_50# N2 a_9280_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X337 a_460_990# P2 a_370_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X338 a_910_50# X a_820_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X339 a_10360_990# P1 a_10270_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X340 a_10000_1690# X a_9910_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X341 a_6670_750# P0 a_6580_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X342 a_9100_1690# X VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X343 VSSA N2 a_10540_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X344 VSSA N1 a_4600_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X345 a_4960_1690# Y a_4870_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X346 Y P2 a_2440_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X347 a_1630_750# P2 a_1540_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X348 a_4060_1690# N1 a_3970_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X349 a_6940_1690# N1 N1 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X350 a_7930_990# P1 a_7840_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X351 a_9640_750# P2 N2 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X352 a_5770_50# Y a_5680_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X353 a_6940_50# N1 a_6850_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X354 a_10670_975# a_10670_975# a_10810_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X355 a_100_990# a_n310_975# a_10_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X356 a_5500_990# P2 a_5410_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X357 a_10_750# a_n310_700# a_n310_700# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X358 a_2890_990# P2 a_2800_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X359 a_7210_750# P2 a_7120_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X360 a_n260_50# a_n310_35# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X361 N2 N2 a_9820_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X362 Z X a_1360_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X363 X X a_1000_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X364 a_4600_1690# Y VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X365 a_2170_750# P1 a_2080_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X366 a_7480_1690# N1 a_7390_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X367 a_8470_990# P2 a_8380_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X368 a_6580_1690# N1 a_6490_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X369 VDDA P1 a_7480_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X370 VSSA a_10670_35# a_11080_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X371 VSSA X a_10360_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X372 P1 LO N1 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X373 a_2440_1690# N1 a_2350_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X374 a_3430_990# P0 a_3340_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X375 VDDA P0 a_7660_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X376 a_1000_990# P1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X377 VSSA Y a_6220_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X378 a_10990_750# a_10670_700# a_10670_700# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X379 VDDA a_n310_700# a_100_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X380 a_7480_50# N1 a_7390_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X381 a_2710_750# P2 a_2620_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X382 VDDA P1 a_8920_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X383 a_8020_1690# Y Z VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X384 a_10090_750# P1 a_10000_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X385 a_7120_1690# N1 a_7030_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X386 a_8110_990# P2 a_8020_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X387 a_3970_990# P2 a_3880_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X388 a_2980_1690# N1 a_2890_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X389 a_2080_1690# N1 P2 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X390 a_1630_50# X a_1540_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X391 VDDA P2 a_2980_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X392 VDDA P1 a_3160_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X393 a_n170_990# a_n310_975# a_n260_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X394 a_4600_50# N1 a_4510_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X395 VDDA P1 a_10540_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X396 a_5230_750# P0 a_5140_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X397 a_8650_990# P2 a_8560_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X398 a_7660_1690# X VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X399 a_3520_1690# N1 a_3430_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X400 VDDA P0 a_4420_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X401 a_6850_50# N1 a_6760_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X402 a_3610_990# P2 a_3520_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X403 a_2620_1690# N1 a_2530_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X404 a_8020_50# N1 a_7930_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X405 a_6490_990# P2 a_6400_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X406 a_5590_990# P2 a_5500_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X407 VDDA a_10670_700# a_11080_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X408 a_8200_1690# Y a_8110_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X409 a_5770_750# P2 a_5680_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X410 Z X a_2080_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X411 a_3340_50# N1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X412 a_3160_1690# N1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X413 X P2 a_640_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X414 a_4150_990# P2 a_4060_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X415 a_6040_1690# N1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X416 a_7030_990# P2 a_6940_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X417 a_5140_1690# Y a_5050_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X418 a_8740_750# P2 a_8650_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X419 a_6130_990# P1 a_6040_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X420 a_n260_1690# a_n310_1640# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X421 VDDA P0 a_6220_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X422 a_1990_990# P2 a_1900_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X423 a_1090_990# P1 a_1000_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X424 a_3700_1690# N1 a_3610_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X425 a_1270_750# P1 a_1180_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X426 a_11080_1690# a_10670_1640# a_10990_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X427 a_5680_1690# Y a_5590_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X428 a_9280_750# P1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X429 N1 P2 a_6580_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X430 a_2710_50# Y a_2620_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X431 a_10990_50# a_10670_35# a_10670_35# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X432 a_3880_50# N1 a_3790_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X433 a_2530_990# P2 a_2440_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X434 a_1540_1690# N2 a_1450_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X435 a_6850_750# P2 a_6760_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X436 a_640_1690# N2 a_550_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X437 a_4240_750# P2 N1 VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X438 VDDA P1 a_1540_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X439 a_9640_990# P1 a_9550_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X440 VDDA P1 a_1720_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X441 a_10_990# a_n310_975# a_n310_975# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X442 a_9820_750# P1 a_9730_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X443 a_7210_990# P2 a_7120_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X444 a_6220_1690# N1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X445 a_7570_50# N1 a_7480_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X446 a_8740_50# N1 a_8650_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X447 a_4780_750# P1 a_4690_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X448 a_2170_990# P2 a_2080_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X449 a_1180_1690# N2 a_1090_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X450 a_9190_1690# X a_9100_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X451 a_10360_50# N2 a_10270_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X452 VSSA X a_3160_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X453 a_4420_50# N1 a_4330_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X454 a_2350_750# P2 a_2260_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X455 P1 LO N1 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X456 a_7750_990# P1 a_7660_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X457 LO N1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X458 a_5140_50# Y a_5050_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1e+11p ps=1.4e+06u w=1e+06u l=500000u
X459 a_5500_50# Y a_5410_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X460 VDDA a_n310_975# a_100_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X461 a_1720_1690# N1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X462 a_10990_990# a_10670_975# a_10670_975# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X463 a_2710_990# P2 a_2620_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X464 X P2 a_10000_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X465 X X a_9640_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X466 P2 N1 a_8020_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X467 a_9280_50# N2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X468 VDDA LO a_280_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X469 a_820_50# X Z VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X470 N2 P2 a_10180_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X471 a_7300_1690# N1 a_7210_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X472 a_1990_50# X a_1900_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X473 a_4690_1690# Y a_4600_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X474 a_10670_35# a_10670_35# a_10810_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X475 a_3250_990# P0 a_3160_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X476 a_2260_1690# N1 a_2170_1690# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X477 LO N1 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X478 a_4960_50# Y VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=1e+11p pd=1.4e+06u as=0p ps=0u w=1e+06u l=500000u
X479 VDDA LO a_10540_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X480 a_7840_750# P2 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X481 P0 P2 a_5140_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X482 a_5680_50# Y P0 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X483 a_10810_750# a_10670_700# a_10720_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X484 a_5410_750# P2 a_5320_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X485 a_n170_50# a_n310_35# a_n260_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X486 a_280_1690# N2 VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X487 a_2800_1690# N1 P2 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X488 a_8650_50# N1 a_8560_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X489 a_9820_50# N2 a_9730_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X490 VDDA a_10670_975# a_11080_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X491 a_10180_1690# X Z VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X492 a_1360_50# X a_1270_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X493 a_8380_750# P2 a_8290_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X494 a_5770_990# P0 a_5680_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X495 Y Y a_2440_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X496 a_11080_50# a_10670_35# a_10990_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X497 a_5950_750# P2 a_5860_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X498 a_3340_750# P1 VDDA VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X499 a_730_990# P2 a_640_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X500 a_5050_750# P0 a_4960_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X501 a_8740_990# P1 a_8650_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X502 a_910_750# P2 a_820_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X503 a_10720_1690# a_10670_1640# VSSA VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X504 a_5050_50# Y a_4960_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X505 a_5320_1690# Y P0 VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X506 a_6220_50# Y a_6130_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X507 a_8920_750# P2 a_8830_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X508 a_6310_990# P1 a_6220_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X509 a_7390_50# N1 a_7300_50# VSSA sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X510 a_3880_750# P2 a_3790_750# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X511 N2 P2 a_1180_990# VDDA sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
.ends

.subckt opamp VDDA VSSA INM INP OUT
Xota_0 VDDA VSSA P1 P2 N2 N1 INP INM X ota
Xbuffer_0 VDDA VSSA P1 P2 N1 N2 buffer_0/in X X INM VSSA INP buffer_0/xp buffer
Xbias_0 VDDA VSSA P1 P2 N2 N1 bias
.ends

