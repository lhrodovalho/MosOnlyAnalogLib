magic
tech sky130A
timestamp 1624070110
<< nwell >>
rect -11635 720 65 1275
<< mvnmos >>
rect -11525 1845 -11475 1945
rect -11435 1845 -11385 1945
rect -11345 1845 -11295 1945
rect -11255 1845 -11205 1945
rect -11165 1845 -11115 1945
rect -11075 1845 -11025 1945
rect -10985 1845 -10935 1945
rect -10895 1845 -10845 1945
rect -10805 1845 -10755 1945
rect -10715 1845 -10665 1945
rect -10625 1845 -10575 1945
rect -10535 1845 -10485 1945
rect -10445 1845 -10395 1945
rect -10355 1845 -10305 1945
rect -10265 1845 -10215 1945
rect -10175 1845 -10125 1945
rect -10085 1845 -10035 1945
rect -9995 1845 -9945 1945
rect -9905 1845 -9855 1945
rect -9815 1845 -9765 1945
rect -9725 1845 -9675 1945
rect -9635 1845 -9585 1945
rect -9545 1845 -9495 1945
rect -9455 1845 -9405 1945
rect -9365 1845 -9315 1945
rect -9275 1845 -9225 1945
rect -9185 1845 -9135 1945
rect -9095 1845 -9045 1945
rect -9005 1845 -8955 1945
rect -8915 1845 -8865 1945
rect -8825 1845 -8775 1945
rect -8735 1845 -8685 1945
rect -8645 1845 -8595 1945
rect -8555 1845 -8505 1945
rect -8465 1845 -8415 1945
rect -8375 1845 -8325 1945
rect -8285 1845 -8235 1945
rect -8195 1845 -8145 1945
rect -8105 1845 -8055 1945
rect -8015 1845 -7965 1945
rect -7925 1845 -7875 1945
rect -7835 1845 -7785 1945
rect -7745 1845 -7695 1945
rect -7655 1845 -7605 1945
rect -7565 1845 -7515 1945
rect -7475 1845 -7425 1945
rect -7385 1845 -7335 1945
rect -7295 1845 -7245 1945
rect -7205 1845 -7155 1945
rect -7115 1845 -7065 1945
rect -7025 1845 -6975 1945
rect -6935 1845 -6885 1945
rect -6845 1845 -6795 1945
rect -6755 1845 -6705 1945
rect -6665 1845 -6615 1945
rect -6575 1845 -6525 1945
rect -6485 1845 -6435 1945
rect -6395 1845 -6345 1945
rect -6305 1845 -6255 1945
rect -6215 1845 -6165 1945
rect -6125 1845 -6075 1945
rect -6035 1845 -5985 1945
rect -5945 1845 -5895 1945
rect -5855 1845 -5805 1945
rect -5765 1845 -5715 1945
rect -5675 1845 -5625 1945
rect -5585 1845 -5535 1945
rect -5495 1845 -5445 1945
rect -5405 1845 -5355 1945
rect -5315 1845 -5265 1945
rect -5225 1845 -5175 1945
rect -5135 1845 -5085 1945
rect -5045 1845 -4995 1945
rect -4955 1845 -4905 1945
rect -4865 1845 -4815 1945
rect -4775 1845 -4725 1945
rect -4685 1845 -4635 1945
rect -4595 1845 -4545 1945
rect -4505 1845 -4455 1945
rect -4415 1845 -4365 1945
rect -4325 1845 -4275 1945
rect -4235 1845 -4185 1945
rect -4145 1845 -4095 1945
rect -4055 1845 -4005 1945
rect -3965 1845 -3915 1945
rect -3875 1845 -3825 1945
rect -3785 1845 -3735 1945
rect -3695 1845 -3645 1945
rect -3605 1845 -3555 1945
rect -3515 1845 -3465 1945
rect -3425 1845 -3375 1945
rect -3335 1845 -3285 1945
rect -3245 1845 -3195 1945
rect -3155 1845 -3105 1945
rect -3065 1845 -3015 1945
rect -2975 1845 -2925 1945
rect -2885 1845 -2835 1945
rect -2795 1845 -2745 1945
rect -2705 1845 -2655 1945
rect -2615 1845 -2565 1945
rect -2525 1845 -2475 1945
rect -2435 1845 -2385 1945
rect -2345 1845 -2295 1945
rect -2255 1845 -2205 1945
rect -2165 1845 -2115 1945
rect -2075 1845 -2025 1945
rect -1985 1845 -1935 1945
rect -1895 1845 -1845 1945
rect -1805 1845 -1755 1945
rect -1715 1845 -1665 1945
rect -1625 1845 -1575 1945
rect -1535 1845 -1485 1945
rect -1445 1845 -1395 1945
rect -1355 1845 -1305 1945
rect -1265 1845 -1215 1945
rect -1175 1845 -1125 1945
rect -1085 1845 -1035 1945
rect -995 1845 -945 1945
rect -905 1845 -855 1945
rect -815 1845 -765 1945
rect -725 1845 -675 1945
rect -635 1845 -585 1945
rect -545 1845 -495 1945
rect -455 1845 -405 1945
rect -365 1845 -315 1945
rect -275 1845 -225 1945
rect -185 1845 -135 1945
rect -95 1845 -45 1945
rect -11525 50 -11475 150
rect -11435 50 -11385 150
rect -11345 50 -11295 150
rect -11255 50 -11205 150
rect -11165 50 -11115 150
rect -11075 50 -11025 150
rect -10985 50 -10935 150
rect -10895 50 -10845 150
rect -10805 50 -10755 150
rect -10715 50 -10665 150
rect -10625 50 -10575 150
rect -10535 50 -10485 150
rect -10445 50 -10395 150
rect -10355 50 -10305 150
rect -10265 50 -10215 150
rect -10175 50 -10125 150
rect -10085 50 -10035 150
rect -9995 50 -9945 150
rect -9905 50 -9855 150
rect -9815 50 -9765 150
rect -9725 50 -9675 150
rect -9635 50 -9585 150
rect -9545 50 -9495 150
rect -9455 50 -9405 150
rect -9365 50 -9315 150
rect -9275 50 -9225 150
rect -9185 50 -9135 150
rect -9095 50 -9045 150
rect -9005 50 -8955 150
rect -8915 50 -8865 150
rect -8825 50 -8775 150
rect -8735 50 -8685 150
rect -8645 50 -8595 150
rect -8555 50 -8505 150
rect -8465 50 -8415 150
rect -8375 50 -8325 150
rect -8285 50 -8235 150
rect -8195 50 -8145 150
rect -8105 50 -8055 150
rect -8015 50 -7965 150
rect -7925 50 -7875 150
rect -7835 50 -7785 150
rect -7745 50 -7695 150
rect -7655 50 -7605 150
rect -7565 50 -7515 150
rect -7475 50 -7425 150
rect -7385 50 -7335 150
rect -7295 50 -7245 150
rect -7205 50 -7155 150
rect -7115 50 -7065 150
rect -7025 50 -6975 150
rect -6935 50 -6885 150
rect -6845 50 -6795 150
rect -6755 50 -6705 150
rect -6665 50 -6615 150
rect -6575 50 -6525 150
rect -6485 50 -6435 150
rect -6395 50 -6345 150
rect -6305 50 -6255 150
rect -6215 50 -6165 150
rect -6125 50 -6075 150
rect -6035 50 -5985 150
rect -5945 50 -5895 150
rect -5855 50 -5805 150
rect -5765 50 -5715 150
rect -5675 50 -5625 150
rect -5585 50 -5535 150
rect -5495 50 -5445 150
rect -5405 50 -5355 150
rect -5315 50 -5265 150
rect -5225 50 -5175 150
rect -5135 50 -5085 150
rect -5045 50 -4995 150
rect -4955 50 -4905 150
rect -4865 50 -4815 150
rect -4775 50 -4725 150
rect -4685 50 -4635 150
rect -4595 50 -4545 150
rect -4505 50 -4455 150
rect -4415 50 -4365 150
rect -4325 50 -4275 150
rect -4235 50 -4185 150
rect -4145 50 -4095 150
rect -4055 50 -4005 150
rect -3965 50 -3915 150
rect -3875 50 -3825 150
rect -3785 50 -3735 150
rect -3695 50 -3645 150
rect -3605 50 -3555 150
rect -3515 50 -3465 150
rect -3425 50 -3375 150
rect -3335 50 -3285 150
rect -3245 50 -3195 150
rect -3155 50 -3105 150
rect -3065 50 -3015 150
rect -2975 50 -2925 150
rect -2885 50 -2835 150
rect -2795 50 -2745 150
rect -2705 50 -2655 150
rect -2615 50 -2565 150
rect -2525 50 -2475 150
rect -2435 50 -2385 150
rect -2345 50 -2295 150
rect -2255 50 -2205 150
rect -2165 50 -2115 150
rect -2075 50 -2025 150
rect -1985 50 -1935 150
rect -1895 50 -1845 150
rect -1805 50 -1755 150
rect -1715 50 -1665 150
rect -1625 50 -1575 150
rect -1535 50 -1485 150
rect -1445 50 -1395 150
rect -1355 50 -1305 150
rect -1265 50 -1215 150
rect -1175 50 -1125 150
rect -1085 50 -1035 150
rect -995 50 -945 150
rect -905 50 -855 150
rect -815 50 -765 150
rect -725 50 -675 150
rect -635 50 -585 150
rect -545 50 -495 150
rect -455 50 -405 150
rect -365 50 -315 150
rect -275 50 -225 150
rect -185 50 -135 150
rect -95 50 -45 150
<< mvpmos >>
rect -11525 1065 -11475 1165
rect -11435 1065 -11385 1165
rect -11345 1065 -11295 1165
rect -11255 1065 -11205 1165
rect -11165 1065 -11115 1165
rect -11075 1065 -11025 1165
rect -10985 1065 -10935 1165
rect -10895 1065 -10845 1165
rect -10805 1065 -10755 1165
rect -10715 1065 -10665 1165
rect -10625 1065 -10575 1165
rect -10535 1065 -10485 1165
rect -10445 1065 -10395 1165
rect -10355 1065 -10305 1165
rect -10265 1065 -10215 1165
rect -10175 1065 -10125 1165
rect -10085 1065 -10035 1165
rect -9995 1065 -9945 1165
rect -9905 1065 -9855 1165
rect -9815 1065 -9765 1165
rect -9725 1065 -9675 1165
rect -9635 1065 -9585 1165
rect -9545 1065 -9495 1165
rect -9455 1065 -9405 1165
rect -9365 1065 -9315 1165
rect -9275 1065 -9225 1165
rect -9185 1065 -9135 1165
rect -9095 1065 -9045 1165
rect -9005 1065 -8955 1165
rect -8915 1065 -8865 1165
rect -8825 1065 -8775 1165
rect -8735 1065 -8685 1165
rect -8645 1065 -8595 1165
rect -8555 1065 -8505 1165
rect -8465 1065 -8415 1165
rect -8375 1065 -8325 1165
rect -8285 1065 -8235 1165
rect -8195 1065 -8145 1165
rect -8105 1065 -8055 1165
rect -8015 1065 -7965 1165
rect -7925 1065 -7875 1165
rect -7835 1065 -7785 1165
rect -7745 1065 -7695 1165
rect -7655 1065 -7605 1165
rect -7565 1065 -7515 1165
rect -7475 1065 -7425 1165
rect -7385 1065 -7335 1165
rect -7295 1065 -7245 1165
rect -7205 1065 -7155 1165
rect -7115 1065 -7065 1165
rect -7025 1065 -6975 1165
rect -6935 1065 -6885 1165
rect -6845 1065 -6795 1165
rect -6755 1065 -6705 1165
rect -6665 1065 -6615 1165
rect -6575 1065 -6525 1165
rect -6485 1065 -6435 1165
rect -6395 1065 -6345 1165
rect -6305 1065 -6255 1165
rect -6215 1065 -6165 1165
rect -6125 1065 -6075 1165
rect -6035 1065 -5985 1165
rect -5945 1065 -5895 1165
rect -5855 1065 -5805 1165
rect -5765 1065 -5715 1165
rect -5675 1065 -5625 1165
rect -5585 1065 -5535 1165
rect -5495 1065 -5445 1165
rect -5405 1065 -5355 1165
rect -5315 1065 -5265 1165
rect -5225 1065 -5175 1165
rect -5135 1065 -5085 1165
rect -5045 1065 -4995 1165
rect -4955 1065 -4905 1165
rect -4865 1065 -4815 1165
rect -4775 1065 -4725 1165
rect -4685 1065 -4635 1165
rect -4595 1065 -4545 1165
rect -4505 1065 -4455 1165
rect -4415 1065 -4365 1165
rect -4325 1065 -4275 1165
rect -4235 1065 -4185 1165
rect -4145 1065 -4095 1165
rect -4055 1065 -4005 1165
rect -3965 1065 -3915 1165
rect -3875 1065 -3825 1165
rect -3785 1065 -3735 1165
rect -3695 1065 -3645 1165
rect -3605 1065 -3555 1165
rect -3515 1065 -3465 1165
rect -3425 1065 -3375 1165
rect -3335 1065 -3285 1165
rect -3245 1065 -3195 1165
rect -3155 1065 -3105 1165
rect -3065 1065 -3015 1165
rect -2975 1065 -2925 1165
rect -2885 1065 -2835 1165
rect -2795 1065 -2745 1165
rect -2705 1065 -2655 1165
rect -2615 1065 -2565 1165
rect -2525 1065 -2475 1165
rect -2435 1065 -2385 1165
rect -2345 1065 -2295 1165
rect -2255 1065 -2205 1165
rect -2165 1065 -2115 1165
rect -2075 1065 -2025 1165
rect -1985 1065 -1935 1165
rect -1895 1065 -1845 1165
rect -1805 1065 -1755 1165
rect -1715 1065 -1665 1165
rect -1625 1065 -1575 1165
rect -1535 1065 -1485 1165
rect -1445 1065 -1395 1165
rect -1355 1065 -1305 1165
rect -1265 1065 -1215 1165
rect -1175 1065 -1125 1165
rect -1085 1065 -1035 1165
rect -995 1065 -945 1165
rect -905 1065 -855 1165
rect -815 1065 -765 1165
rect -725 1065 -675 1165
rect -635 1065 -585 1165
rect -545 1065 -495 1165
rect -455 1065 -405 1165
rect -365 1065 -315 1165
rect -275 1065 -225 1165
rect -185 1065 -135 1165
rect -95 1065 -45 1165
rect -11525 830 -11475 930
rect -11435 830 -11385 930
rect -11345 830 -11295 930
rect -11255 830 -11205 930
rect -11165 830 -11115 930
rect -11075 830 -11025 930
rect -10985 830 -10935 930
rect -10895 830 -10845 930
rect -10805 830 -10755 930
rect -10715 830 -10665 930
rect -10625 830 -10575 930
rect -10535 830 -10485 930
rect -10445 830 -10395 930
rect -10355 830 -10305 930
rect -10265 830 -10215 930
rect -10175 830 -10125 930
rect -10085 830 -10035 930
rect -9995 830 -9945 930
rect -9905 830 -9855 930
rect -9815 830 -9765 930
rect -9725 830 -9675 930
rect -9635 830 -9585 930
rect -9545 830 -9495 930
rect -9455 830 -9405 930
rect -9365 830 -9315 930
rect -9275 830 -9225 930
rect -9185 830 -9135 930
rect -9095 830 -9045 930
rect -9005 830 -8955 930
rect -8915 830 -8865 930
rect -8825 830 -8775 930
rect -8735 830 -8685 930
rect -8645 830 -8595 930
rect -8555 830 -8505 930
rect -8465 830 -8415 930
rect -8375 830 -8325 930
rect -8285 830 -8235 930
rect -8195 830 -8145 930
rect -8105 830 -8055 930
rect -8015 830 -7965 930
rect -7925 830 -7875 930
rect -7835 830 -7785 930
rect -7745 830 -7695 930
rect -7655 830 -7605 930
rect -7565 830 -7515 930
rect -7475 830 -7425 930
rect -7385 830 -7335 930
rect -7295 830 -7245 930
rect -7205 830 -7155 930
rect -7115 830 -7065 930
rect -7025 830 -6975 930
rect -6935 830 -6885 930
rect -6845 830 -6795 930
rect -6755 830 -6705 930
rect -6665 830 -6615 930
rect -6575 830 -6525 930
rect -6485 830 -6435 930
rect -6395 830 -6345 930
rect -6305 830 -6255 930
rect -6215 830 -6165 930
rect -6125 830 -6075 930
rect -6035 830 -5985 930
rect -5945 830 -5895 930
rect -5855 830 -5805 930
rect -5765 830 -5715 930
rect -5675 830 -5625 930
rect -5585 830 -5535 930
rect -5495 830 -5445 930
rect -5405 830 -5355 930
rect -5315 830 -5265 930
rect -5225 830 -5175 930
rect -5135 830 -5085 930
rect -5045 830 -4995 930
rect -4955 830 -4905 930
rect -4865 830 -4815 930
rect -4775 830 -4725 930
rect -4685 830 -4635 930
rect -4595 830 -4545 930
rect -4505 830 -4455 930
rect -4415 830 -4365 930
rect -4325 830 -4275 930
rect -4235 830 -4185 930
rect -4145 830 -4095 930
rect -4055 830 -4005 930
rect -3965 830 -3915 930
rect -3875 830 -3825 930
rect -3785 830 -3735 930
rect -3695 830 -3645 930
rect -3605 830 -3555 930
rect -3515 830 -3465 930
rect -3425 830 -3375 930
rect -3335 830 -3285 930
rect -3245 830 -3195 930
rect -3155 830 -3105 930
rect -3065 830 -3015 930
rect -2975 830 -2925 930
rect -2885 830 -2835 930
rect -2795 830 -2745 930
rect -2705 830 -2655 930
rect -2615 830 -2565 930
rect -2525 830 -2475 930
rect -2435 830 -2385 930
rect -2345 830 -2295 930
rect -2255 830 -2205 930
rect -2165 830 -2115 930
rect -2075 830 -2025 930
rect -1985 830 -1935 930
rect -1895 830 -1845 930
rect -1805 830 -1755 930
rect -1715 830 -1665 930
rect -1625 830 -1575 930
rect -1535 830 -1485 930
rect -1445 830 -1395 930
rect -1355 830 -1305 930
rect -1265 830 -1215 930
rect -1175 830 -1125 930
rect -1085 830 -1035 930
rect -995 830 -945 930
rect -905 830 -855 930
rect -815 830 -765 930
rect -725 830 -675 930
rect -635 830 -585 930
rect -545 830 -495 930
rect -455 830 -405 930
rect -365 830 -315 930
rect -275 830 -225 930
rect -185 830 -135 930
rect -95 830 -45 930
<< mvndiff >>
rect -11565 1935 -11525 1945
rect -11565 1855 -11555 1935
rect -11535 1855 -11525 1935
rect -11565 1845 -11525 1855
rect -11475 1935 -11435 1945
rect -11475 1855 -11465 1935
rect -11445 1855 -11435 1935
rect -11475 1845 -11435 1855
rect -11385 1935 -11345 1945
rect -11385 1855 -11375 1935
rect -11355 1855 -11345 1935
rect -11385 1845 -11345 1855
rect -11295 1935 -11255 1945
rect -11295 1855 -11285 1935
rect -11265 1855 -11255 1935
rect -11295 1845 -11255 1855
rect -11205 1935 -11165 1945
rect -11205 1855 -11195 1935
rect -11175 1855 -11165 1935
rect -11205 1845 -11165 1855
rect -11115 1935 -11075 1945
rect -11115 1855 -11105 1935
rect -11085 1855 -11075 1935
rect -11115 1845 -11075 1855
rect -11025 1935 -10985 1945
rect -11025 1855 -11015 1935
rect -10995 1855 -10985 1935
rect -11025 1845 -10985 1855
rect -10935 1935 -10895 1945
rect -10935 1855 -10925 1935
rect -10905 1855 -10895 1935
rect -10935 1845 -10895 1855
rect -10845 1935 -10805 1945
rect -10845 1855 -10835 1935
rect -10815 1855 -10805 1935
rect -10845 1845 -10805 1855
rect -10755 1935 -10715 1945
rect -10755 1855 -10745 1935
rect -10725 1855 -10715 1935
rect -10755 1845 -10715 1855
rect -10665 1935 -10625 1945
rect -10665 1855 -10655 1935
rect -10635 1855 -10625 1935
rect -10665 1845 -10625 1855
rect -10575 1935 -10535 1945
rect -10575 1855 -10565 1935
rect -10545 1855 -10535 1935
rect -10575 1845 -10535 1855
rect -10485 1935 -10445 1945
rect -10485 1855 -10475 1935
rect -10455 1855 -10445 1935
rect -10485 1845 -10445 1855
rect -10395 1935 -10355 1945
rect -10395 1855 -10385 1935
rect -10365 1855 -10355 1935
rect -10395 1845 -10355 1855
rect -10305 1935 -10265 1945
rect -10305 1855 -10295 1935
rect -10275 1855 -10265 1935
rect -10305 1845 -10265 1855
rect -10215 1935 -10175 1945
rect -10215 1855 -10205 1935
rect -10185 1855 -10175 1935
rect -10215 1845 -10175 1855
rect -10125 1935 -10085 1945
rect -10125 1855 -10115 1935
rect -10095 1855 -10085 1935
rect -10125 1845 -10085 1855
rect -10035 1935 -9995 1945
rect -10035 1855 -10025 1935
rect -10005 1855 -9995 1935
rect -10035 1845 -9995 1855
rect -9945 1935 -9905 1945
rect -9945 1855 -9935 1935
rect -9915 1855 -9905 1935
rect -9945 1845 -9905 1855
rect -9855 1935 -9815 1945
rect -9855 1855 -9845 1935
rect -9825 1855 -9815 1935
rect -9855 1845 -9815 1855
rect -9765 1935 -9725 1945
rect -9765 1855 -9755 1935
rect -9735 1855 -9725 1935
rect -9765 1845 -9725 1855
rect -9675 1935 -9635 1945
rect -9675 1855 -9665 1935
rect -9645 1855 -9635 1935
rect -9675 1845 -9635 1855
rect -9585 1935 -9545 1945
rect -9585 1855 -9575 1935
rect -9555 1855 -9545 1935
rect -9585 1845 -9545 1855
rect -9495 1935 -9455 1945
rect -9495 1855 -9485 1935
rect -9465 1855 -9455 1935
rect -9495 1845 -9455 1855
rect -9405 1935 -9365 1945
rect -9405 1855 -9395 1935
rect -9375 1855 -9365 1935
rect -9405 1845 -9365 1855
rect -9315 1935 -9275 1945
rect -9315 1855 -9305 1935
rect -9285 1855 -9275 1935
rect -9315 1845 -9275 1855
rect -9225 1935 -9185 1945
rect -9225 1855 -9215 1935
rect -9195 1855 -9185 1935
rect -9225 1845 -9185 1855
rect -9135 1935 -9095 1945
rect -9135 1855 -9125 1935
rect -9105 1855 -9095 1935
rect -9135 1845 -9095 1855
rect -9045 1935 -9005 1945
rect -9045 1855 -9035 1935
rect -9015 1855 -9005 1935
rect -9045 1845 -9005 1855
rect -8955 1935 -8915 1945
rect -8955 1855 -8945 1935
rect -8925 1855 -8915 1935
rect -8955 1845 -8915 1855
rect -8865 1935 -8825 1945
rect -8865 1855 -8855 1935
rect -8835 1855 -8825 1935
rect -8865 1845 -8825 1855
rect -8775 1935 -8735 1945
rect -8775 1855 -8765 1935
rect -8745 1855 -8735 1935
rect -8775 1845 -8735 1855
rect -8685 1935 -8645 1945
rect -8685 1855 -8675 1935
rect -8655 1855 -8645 1935
rect -8685 1845 -8645 1855
rect -8595 1935 -8555 1945
rect -8595 1855 -8585 1935
rect -8565 1855 -8555 1935
rect -8595 1845 -8555 1855
rect -8505 1935 -8465 1945
rect -8505 1855 -8495 1935
rect -8475 1855 -8465 1935
rect -8505 1845 -8465 1855
rect -8415 1935 -8375 1945
rect -8415 1855 -8405 1935
rect -8385 1855 -8375 1935
rect -8415 1845 -8375 1855
rect -8325 1935 -8285 1945
rect -8325 1855 -8315 1935
rect -8295 1855 -8285 1935
rect -8325 1845 -8285 1855
rect -8235 1935 -8195 1945
rect -8235 1855 -8225 1935
rect -8205 1855 -8195 1935
rect -8235 1845 -8195 1855
rect -8145 1935 -8105 1945
rect -8145 1855 -8135 1935
rect -8115 1855 -8105 1935
rect -8145 1845 -8105 1855
rect -8055 1935 -8015 1945
rect -8055 1855 -8045 1935
rect -8025 1855 -8015 1935
rect -8055 1845 -8015 1855
rect -7965 1935 -7925 1945
rect -7965 1855 -7955 1935
rect -7935 1855 -7925 1935
rect -7965 1845 -7925 1855
rect -7875 1935 -7835 1945
rect -7875 1855 -7865 1935
rect -7845 1855 -7835 1935
rect -7875 1845 -7835 1855
rect -7785 1935 -7745 1945
rect -7785 1855 -7775 1935
rect -7755 1855 -7745 1935
rect -7785 1845 -7745 1855
rect -7695 1935 -7655 1945
rect -7695 1855 -7685 1935
rect -7665 1855 -7655 1935
rect -7695 1845 -7655 1855
rect -7605 1935 -7565 1945
rect -7605 1855 -7595 1935
rect -7575 1855 -7565 1935
rect -7605 1845 -7565 1855
rect -7515 1935 -7475 1945
rect -7515 1855 -7505 1935
rect -7485 1855 -7475 1935
rect -7515 1845 -7475 1855
rect -7425 1935 -7385 1945
rect -7425 1855 -7415 1935
rect -7395 1855 -7385 1935
rect -7425 1845 -7385 1855
rect -7335 1935 -7295 1945
rect -7335 1855 -7325 1935
rect -7305 1855 -7295 1935
rect -7335 1845 -7295 1855
rect -7245 1935 -7205 1945
rect -7245 1855 -7235 1935
rect -7215 1855 -7205 1935
rect -7245 1845 -7205 1855
rect -7155 1935 -7115 1945
rect -7155 1855 -7145 1935
rect -7125 1855 -7115 1935
rect -7155 1845 -7115 1855
rect -7065 1935 -7025 1945
rect -7065 1855 -7055 1935
rect -7035 1855 -7025 1935
rect -7065 1845 -7025 1855
rect -6975 1935 -6935 1945
rect -6975 1855 -6965 1935
rect -6945 1855 -6935 1935
rect -6975 1845 -6935 1855
rect -6885 1935 -6845 1945
rect -6885 1855 -6875 1935
rect -6855 1855 -6845 1935
rect -6885 1845 -6845 1855
rect -6795 1935 -6755 1945
rect -6795 1855 -6785 1935
rect -6765 1855 -6755 1935
rect -6795 1845 -6755 1855
rect -6705 1935 -6665 1945
rect -6705 1855 -6695 1935
rect -6675 1855 -6665 1935
rect -6705 1845 -6665 1855
rect -6615 1935 -6575 1945
rect -6615 1855 -6605 1935
rect -6585 1855 -6575 1935
rect -6615 1845 -6575 1855
rect -6525 1935 -6485 1945
rect -6525 1855 -6515 1935
rect -6495 1855 -6485 1935
rect -6525 1845 -6485 1855
rect -6435 1935 -6395 1945
rect -6435 1855 -6425 1935
rect -6405 1855 -6395 1935
rect -6435 1845 -6395 1855
rect -6345 1935 -6305 1945
rect -6345 1855 -6335 1935
rect -6315 1855 -6305 1935
rect -6345 1845 -6305 1855
rect -6255 1935 -6215 1945
rect -6255 1855 -6245 1935
rect -6225 1855 -6215 1935
rect -6255 1845 -6215 1855
rect -6165 1935 -6125 1945
rect -6165 1855 -6155 1935
rect -6135 1855 -6125 1935
rect -6165 1845 -6125 1855
rect -6075 1935 -6035 1945
rect -6075 1855 -6065 1935
rect -6045 1855 -6035 1935
rect -6075 1845 -6035 1855
rect -5985 1935 -5945 1945
rect -5985 1855 -5975 1935
rect -5955 1855 -5945 1935
rect -5985 1845 -5945 1855
rect -5895 1935 -5855 1945
rect -5895 1855 -5885 1935
rect -5865 1855 -5855 1935
rect -5895 1845 -5855 1855
rect -5805 1935 -5765 1945
rect -5805 1855 -5795 1935
rect -5775 1855 -5765 1935
rect -5805 1845 -5765 1855
rect -5715 1935 -5675 1945
rect -5715 1855 -5705 1935
rect -5685 1855 -5675 1935
rect -5715 1845 -5675 1855
rect -5625 1935 -5585 1945
rect -5625 1855 -5615 1935
rect -5595 1855 -5585 1935
rect -5625 1845 -5585 1855
rect -5535 1935 -5495 1945
rect -5535 1855 -5525 1935
rect -5505 1855 -5495 1935
rect -5535 1845 -5495 1855
rect -5445 1935 -5405 1945
rect -5445 1855 -5435 1935
rect -5415 1855 -5405 1935
rect -5445 1845 -5405 1855
rect -5355 1935 -5315 1945
rect -5355 1855 -5345 1935
rect -5325 1855 -5315 1935
rect -5355 1845 -5315 1855
rect -5265 1935 -5225 1945
rect -5265 1855 -5255 1935
rect -5235 1855 -5225 1935
rect -5265 1845 -5225 1855
rect -5175 1935 -5135 1945
rect -5175 1855 -5165 1935
rect -5145 1855 -5135 1935
rect -5175 1845 -5135 1855
rect -5085 1935 -5045 1945
rect -5085 1855 -5075 1935
rect -5055 1855 -5045 1935
rect -5085 1845 -5045 1855
rect -4995 1935 -4955 1945
rect -4995 1855 -4985 1935
rect -4965 1855 -4955 1935
rect -4995 1845 -4955 1855
rect -4905 1935 -4865 1945
rect -4905 1855 -4895 1935
rect -4875 1855 -4865 1935
rect -4905 1845 -4865 1855
rect -4815 1935 -4775 1945
rect -4815 1855 -4805 1935
rect -4785 1855 -4775 1935
rect -4815 1845 -4775 1855
rect -4725 1935 -4685 1945
rect -4725 1855 -4715 1935
rect -4695 1855 -4685 1935
rect -4725 1845 -4685 1855
rect -4635 1935 -4595 1945
rect -4635 1855 -4625 1935
rect -4605 1855 -4595 1935
rect -4635 1845 -4595 1855
rect -4545 1935 -4505 1945
rect -4545 1855 -4535 1935
rect -4515 1855 -4505 1935
rect -4545 1845 -4505 1855
rect -4455 1935 -4415 1945
rect -4455 1855 -4445 1935
rect -4425 1855 -4415 1935
rect -4455 1845 -4415 1855
rect -4365 1935 -4325 1945
rect -4365 1855 -4355 1935
rect -4335 1855 -4325 1935
rect -4365 1845 -4325 1855
rect -4275 1935 -4235 1945
rect -4275 1855 -4265 1935
rect -4245 1855 -4235 1935
rect -4275 1845 -4235 1855
rect -4185 1935 -4145 1945
rect -4185 1855 -4175 1935
rect -4155 1855 -4145 1935
rect -4185 1845 -4145 1855
rect -4095 1935 -4055 1945
rect -4095 1855 -4085 1935
rect -4065 1855 -4055 1935
rect -4095 1845 -4055 1855
rect -4005 1935 -3965 1945
rect -4005 1855 -3995 1935
rect -3975 1855 -3965 1935
rect -4005 1845 -3965 1855
rect -3915 1935 -3875 1945
rect -3915 1855 -3905 1935
rect -3885 1855 -3875 1935
rect -3915 1845 -3875 1855
rect -3825 1935 -3785 1945
rect -3825 1855 -3815 1935
rect -3795 1855 -3785 1935
rect -3825 1845 -3785 1855
rect -3735 1935 -3695 1945
rect -3735 1855 -3725 1935
rect -3705 1855 -3695 1935
rect -3735 1845 -3695 1855
rect -3645 1935 -3605 1945
rect -3645 1855 -3635 1935
rect -3615 1855 -3605 1935
rect -3645 1845 -3605 1855
rect -3555 1935 -3515 1945
rect -3555 1855 -3545 1935
rect -3525 1855 -3515 1935
rect -3555 1845 -3515 1855
rect -3465 1935 -3425 1945
rect -3465 1855 -3455 1935
rect -3435 1855 -3425 1935
rect -3465 1845 -3425 1855
rect -3375 1935 -3335 1945
rect -3375 1855 -3365 1935
rect -3345 1855 -3335 1935
rect -3375 1845 -3335 1855
rect -3285 1935 -3245 1945
rect -3285 1855 -3275 1935
rect -3255 1855 -3245 1935
rect -3285 1845 -3245 1855
rect -3195 1935 -3155 1945
rect -3195 1855 -3185 1935
rect -3165 1855 -3155 1935
rect -3195 1845 -3155 1855
rect -3105 1935 -3065 1945
rect -3105 1855 -3095 1935
rect -3075 1855 -3065 1935
rect -3105 1845 -3065 1855
rect -3015 1935 -2975 1945
rect -3015 1855 -3005 1935
rect -2985 1855 -2975 1935
rect -3015 1845 -2975 1855
rect -2925 1935 -2885 1945
rect -2925 1855 -2915 1935
rect -2895 1855 -2885 1935
rect -2925 1845 -2885 1855
rect -2835 1935 -2795 1945
rect -2835 1855 -2825 1935
rect -2805 1855 -2795 1935
rect -2835 1845 -2795 1855
rect -2745 1935 -2705 1945
rect -2745 1855 -2735 1935
rect -2715 1855 -2705 1935
rect -2745 1845 -2705 1855
rect -2655 1935 -2615 1945
rect -2655 1855 -2645 1935
rect -2625 1855 -2615 1935
rect -2655 1845 -2615 1855
rect -2565 1935 -2525 1945
rect -2565 1855 -2555 1935
rect -2535 1855 -2525 1935
rect -2565 1845 -2525 1855
rect -2475 1935 -2435 1945
rect -2475 1855 -2465 1935
rect -2445 1855 -2435 1935
rect -2475 1845 -2435 1855
rect -2385 1935 -2345 1945
rect -2385 1855 -2375 1935
rect -2355 1855 -2345 1935
rect -2385 1845 -2345 1855
rect -2295 1935 -2255 1945
rect -2295 1855 -2285 1935
rect -2265 1855 -2255 1935
rect -2295 1845 -2255 1855
rect -2205 1935 -2165 1945
rect -2205 1855 -2195 1935
rect -2175 1855 -2165 1935
rect -2205 1845 -2165 1855
rect -2115 1935 -2075 1945
rect -2115 1855 -2105 1935
rect -2085 1855 -2075 1935
rect -2115 1845 -2075 1855
rect -2025 1935 -1985 1945
rect -2025 1855 -2015 1935
rect -1995 1855 -1985 1935
rect -2025 1845 -1985 1855
rect -1935 1935 -1895 1945
rect -1935 1855 -1925 1935
rect -1905 1855 -1895 1935
rect -1935 1845 -1895 1855
rect -1845 1935 -1805 1945
rect -1845 1855 -1835 1935
rect -1815 1855 -1805 1935
rect -1845 1845 -1805 1855
rect -1755 1935 -1715 1945
rect -1755 1855 -1745 1935
rect -1725 1855 -1715 1935
rect -1755 1845 -1715 1855
rect -1665 1935 -1625 1945
rect -1665 1855 -1655 1935
rect -1635 1855 -1625 1935
rect -1665 1845 -1625 1855
rect -1575 1935 -1535 1945
rect -1575 1855 -1565 1935
rect -1545 1855 -1535 1935
rect -1575 1845 -1535 1855
rect -1485 1935 -1445 1945
rect -1485 1855 -1475 1935
rect -1455 1855 -1445 1935
rect -1485 1845 -1445 1855
rect -1395 1935 -1355 1945
rect -1395 1855 -1385 1935
rect -1365 1855 -1355 1935
rect -1395 1845 -1355 1855
rect -1305 1935 -1265 1945
rect -1305 1855 -1295 1935
rect -1275 1855 -1265 1935
rect -1305 1845 -1265 1855
rect -1215 1935 -1175 1945
rect -1215 1855 -1205 1935
rect -1185 1855 -1175 1935
rect -1215 1845 -1175 1855
rect -1125 1935 -1085 1945
rect -1125 1855 -1115 1935
rect -1095 1855 -1085 1935
rect -1125 1845 -1085 1855
rect -1035 1935 -995 1945
rect -1035 1855 -1025 1935
rect -1005 1855 -995 1935
rect -1035 1845 -995 1855
rect -945 1935 -905 1945
rect -945 1855 -935 1935
rect -915 1855 -905 1935
rect -945 1845 -905 1855
rect -855 1935 -815 1945
rect -855 1855 -845 1935
rect -825 1855 -815 1935
rect -855 1845 -815 1855
rect -765 1935 -725 1945
rect -765 1855 -755 1935
rect -735 1855 -725 1935
rect -765 1845 -725 1855
rect -675 1935 -635 1945
rect -675 1855 -665 1935
rect -645 1855 -635 1935
rect -675 1845 -635 1855
rect -585 1935 -545 1945
rect -585 1855 -575 1935
rect -555 1855 -545 1935
rect -585 1845 -545 1855
rect -495 1935 -455 1945
rect -495 1855 -485 1935
rect -465 1855 -455 1935
rect -495 1845 -455 1855
rect -405 1935 -365 1945
rect -405 1855 -395 1935
rect -375 1855 -365 1935
rect -405 1845 -365 1855
rect -315 1935 -275 1945
rect -315 1855 -305 1935
rect -285 1855 -275 1935
rect -315 1845 -275 1855
rect -225 1935 -185 1945
rect -225 1855 -215 1935
rect -195 1855 -185 1935
rect -225 1845 -185 1855
rect -135 1935 -95 1945
rect -135 1855 -125 1935
rect -105 1855 -95 1935
rect -135 1845 -95 1855
rect -45 1935 -5 1945
rect -45 1855 -35 1935
rect -15 1855 -5 1935
rect -45 1845 -5 1855
rect -11565 140 -11525 150
rect -11565 60 -11555 140
rect -11535 60 -11525 140
rect -11565 50 -11525 60
rect -11475 140 -11435 150
rect -11475 60 -11465 140
rect -11445 60 -11435 140
rect -11475 50 -11435 60
rect -11385 140 -11345 150
rect -11385 60 -11375 140
rect -11355 60 -11345 140
rect -11385 50 -11345 60
rect -11295 140 -11255 150
rect -11295 60 -11285 140
rect -11265 60 -11255 140
rect -11295 50 -11255 60
rect -11205 140 -11165 150
rect -11205 60 -11195 140
rect -11175 60 -11165 140
rect -11205 50 -11165 60
rect -11115 140 -11075 150
rect -11115 60 -11105 140
rect -11085 60 -11075 140
rect -11115 50 -11075 60
rect -11025 140 -10985 150
rect -11025 60 -11015 140
rect -10995 60 -10985 140
rect -11025 50 -10985 60
rect -10935 140 -10895 150
rect -10935 60 -10925 140
rect -10905 60 -10895 140
rect -10935 50 -10895 60
rect -10845 140 -10805 150
rect -10845 60 -10835 140
rect -10815 60 -10805 140
rect -10845 50 -10805 60
rect -10755 140 -10715 150
rect -10755 60 -10745 140
rect -10725 60 -10715 140
rect -10755 50 -10715 60
rect -10665 140 -10625 150
rect -10665 60 -10655 140
rect -10635 60 -10625 140
rect -10665 50 -10625 60
rect -10575 140 -10535 150
rect -10575 60 -10565 140
rect -10545 60 -10535 140
rect -10575 50 -10535 60
rect -10485 140 -10445 150
rect -10485 60 -10475 140
rect -10455 60 -10445 140
rect -10485 50 -10445 60
rect -10395 140 -10355 150
rect -10395 60 -10385 140
rect -10365 60 -10355 140
rect -10395 50 -10355 60
rect -10305 140 -10265 150
rect -10305 60 -10295 140
rect -10275 60 -10265 140
rect -10305 50 -10265 60
rect -10215 140 -10175 150
rect -10215 60 -10205 140
rect -10185 60 -10175 140
rect -10215 50 -10175 60
rect -10125 140 -10085 150
rect -10125 60 -10115 140
rect -10095 60 -10085 140
rect -10125 50 -10085 60
rect -10035 140 -9995 150
rect -10035 60 -10025 140
rect -10005 60 -9995 140
rect -10035 50 -9995 60
rect -9945 140 -9905 150
rect -9945 60 -9935 140
rect -9915 60 -9905 140
rect -9945 50 -9905 60
rect -9855 140 -9815 150
rect -9855 60 -9845 140
rect -9825 60 -9815 140
rect -9855 50 -9815 60
rect -9765 140 -9725 150
rect -9765 60 -9755 140
rect -9735 60 -9725 140
rect -9765 50 -9725 60
rect -9675 140 -9635 150
rect -9675 60 -9665 140
rect -9645 60 -9635 140
rect -9675 50 -9635 60
rect -9585 140 -9545 150
rect -9585 60 -9575 140
rect -9555 60 -9545 140
rect -9585 50 -9545 60
rect -9495 140 -9455 150
rect -9495 60 -9485 140
rect -9465 60 -9455 140
rect -9495 50 -9455 60
rect -9405 140 -9365 150
rect -9405 60 -9395 140
rect -9375 60 -9365 140
rect -9405 50 -9365 60
rect -9315 140 -9275 150
rect -9315 60 -9305 140
rect -9285 60 -9275 140
rect -9315 50 -9275 60
rect -9225 140 -9185 150
rect -9225 60 -9215 140
rect -9195 60 -9185 140
rect -9225 50 -9185 60
rect -9135 140 -9095 150
rect -9135 60 -9125 140
rect -9105 60 -9095 140
rect -9135 50 -9095 60
rect -9045 140 -9005 150
rect -9045 60 -9035 140
rect -9015 60 -9005 140
rect -9045 50 -9005 60
rect -8955 140 -8915 150
rect -8955 60 -8945 140
rect -8925 60 -8915 140
rect -8955 50 -8915 60
rect -8865 140 -8825 150
rect -8865 60 -8855 140
rect -8835 60 -8825 140
rect -8865 50 -8825 60
rect -8775 140 -8735 150
rect -8775 60 -8765 140
rect -8745 60 -8735 140
rect -8775 50 -8735 60
rect -8685 140 -8645 150
rect -8685 60 -8675 140
rect -8655 60 -8645 140
rect -8685 50 -8645 60
rect -8595 140 -8555 150
rect -8595 60 -8585 140
rect -8565 60 -8555 140
rect -8595 50 -8555 60
rect -8505 140 -8465 150
rect -8505 60 -8495 140
rect -8475 60 -8465 140
rect -8505 50 -8465 60
rect -8415 140 -8375 150
rect -8415 60 -8405 140
rect -8385 60 -8375 140
rect -8415 50 -8375 60
rect -8325 140 -8285 150
rect -8325 60 -8315 140
rect -8295 60 -8285 140
rect -8325 50 -8285 60
rect -8235 140 -8195 150
rect -8235 60 -8225 140
rect -8205 60 -8195 140
rect -8235 50 -8195 60
rect -8145 140 -8105 150
rect -8145 60 -8135 140
rect -8115 60 -8105 140
rect -8145 50 -8105 60
rect -8055 140 -8015 150
rect -8055 60 -8045 140
rect -8025 60 -8015 140
rect -8055 50 -8015 60
rect -7965 140 -7925 150
rect -7965 60 -7955 140
rect -7935 60 -7925 140
rect -7965 50 -7925 60
rect -7875 140 -7835 150
rect -7875 60 -7865 140
rect -7845 60 -7835 140
rect -7875 50 -7835 60
rect -7785 140 -7745 150
rect -7785 60 -7775 140
rect -7755 60 -7745 140
rect -7785 50 -7745 60
rect -7695 140 -7655 150
rect -7695 60 -7685 140
rect -7665 60 -7655 140
rect -7695 50 -7655 60
rect -7605 140 -7565 150
rect -7605 60 -7595 140
rect -7575 60 -7565 140
rect -7605 50 -7565 60
rect -7515 140 -7475 150
rect -7515 60 -7505 140
rect -7485 60 -7475 140
rect -7515 50 -7475 60
rect -7425 140 -7385 150
rect -7425 60 -7415 140
rect -7395 60 -7385 140
rect -7425 50 -7385 60
rect -7335 140 -7295 150
rect -7335 60 -7325 140
rect -7305 60 -7295 140
rect -7335 50 -7295 60
rect -7245 140 -7205 150
rect -7245 60 -7235 140
rect -7215 60 -7205 140
rect -7245 50 -7205 60
rect -7155 140 -7115 150
rect -7155 60 -7145 140
rect -7125 60 -7115 140
rect -7155 50 -7115 60
rect -7065 140 -7025 150
rect -7065 60 -7055 140
rect -7035 60 -7025 140
rect -7065 50 -7025 60
rect -6975 140 -6935 150
rect -6975 60 -6965 140
rect -6945 60 -6935 140
rect -6975 50 -6935 60
rect -6885 140 -6845 150
rect -6885 60 -6875 140
rect -6855 60 -6845 140
rect -6885 50 -6845 60
rect -6795 140 -6755 150
rect -6795 60 -6785 140
rect -6765 60 -6755 140
rect -6795 50 -6755 60
rect -6705 140 -6665 150
rect -6705 60 -6695 140
rect -6675 60 -6665 140
rect -6705 50 -6665 60
rect -6615 140 -6575 150
rect -6615 60 -6605 140
rect -6585 60 -6575 140
rect -6615 50 -6575 60
rect -6525 140 -6485 150
rect -6525 60 -6515 140
rect -6495 60 -6485 140
rect -6525 50 -6485 60
rect -6435 140 -6395 150
rect -6435 60 -6425 140
rect -6405 60 -6395 140
rect -6435 50 -6395 60
rect -6345 140 -6305 150
rect -6345 60 -6335 140
rect -6315 60 -6305 140
rect -6345 50 -6305 60
rect -6255 140 -6215 150
rect -6255 60 -6245 140
rect -6225 60 -6215 140
rect -6255 50 -6215 60
rect -6165 140 -6125 150
rect -6165 60 -6155 140
rect -6135 60 -6125 140
rect -6165 50 -6125 60
rect -6075 140 -6035 150
rect -6075 60 -6065 140
rect -6045 60 -6035 140
rect -6075 50 -6035 60
rect -5985 140 -5945 150
rect -5985 60 -5975 140
rect -5955 60 -5945 140
rect -5985 50 -5945 60
rect -5895 140 -5855 150
rect -5895 60 -5885 140
rect -5865 60 -5855 140
rect -5895 50 -5855 60
rect -5805 140 -5765 150
rect -5805 60 -5795 140
rect -5775 60 -5765 140
rect -5805 50 -5765 60
rect -5715 140 -5675 150
rect -5715 60 -5705 140
rect -5685 60 -5675 140
rect -5715 50 -5675 60
rect -5625 140 -5585 150
rect -5625 60 -5615 140
rect -5595 60 -5585 140
rect -5625 50 -5585 60
rect -5535 140 -5495 150
rect -5535 60 -5525 140
rect -5505 60 -5495 140
rect -5535 50 -5495 60
rect -5445 140 -5405 150
rect -5445 60 -5435 140
rect -5415 60 -5405 140
rect -5445 50 -5405 60
rect -5355 140 -5315 150
rect -5355 60 -5345 140
rect -5325 60 -5315 140
rect -5355 50 -5315 60
rect -5265 140 -5225 150
rect -5265 60 -5255 140
rect -5235 60 -5225 140
rect -5265 50 -5225 60
rect -5175 140 -5135 150
rect -5175 60 -5165 140
rect -5145 60 -5135 140
rect -5175 50 -5135 60
rect -5085 140 -5045 150
rect -5085 60 -5075 140
rect -5055 60 -5045 140
rect -5085 50 -5045 60
rect -4995 140 -4955 150
rect -4995 60 -4985 140
rect -4965 60 -4955 140
rect -4995 50 -4955 60
rect -4905 140 -4865 150
rect -4905 60 -4895 140
rect -4875 60 -4865 140
rect -4905 50 -4865 60
rect -4815 140 -4775 150
rect -4815 60 -4805 140
rect -4785 60 -4775 140
rect -4815 50 -4775 60
rect -4725 140 -4685 150
rect -4725 60 -4715 140
rect -4695 60 -4685 140
rect -4725 50 -4685 60
rect -4635 140 -4595 150
rect -4635 60 -4625 140
rect -4605 60 -4595 140
rect -4635 50 -4595 60
rect -4545 140 -4505 150
rect -4545 60 -4535 140
rect -4515 60 -4505 140
rect -4545 50 -4505 60
rect -4455 140 -4415 150
rect -4455 60 -4445 140
rect -4425 60 -4415 140
rect -4455 50 -4415 60
rect -4365 140 -4325 150
rect -4365 60 -4355 140
rect -4335 60 -4325 140
rect -4365 50 -4325 60
rect -4275 140 -4235 150
rect -4275 60 -4265 140
rect -4245 60 -4235 140
rect -4275 50 -4235 60
rect -4185 140 -4145 150
rect -4185 60 -4175 140
rect -4155 60 -4145 140
rect -4185 50 -4145 60
rect -4095 140 -4055 150
rect -4095 60 -4085 140
rect -4065 60 -4055 140
rect -4095 50 -4055 60
rect -4005 140 -3965 150
rect -4005 60 -3995 140
rect -3975 60 -3965 140
rect -4005 50 -3965 60
rect -3915 140 -3875 150
rect -3915 60 -3905 140
rect -3885 60 -3875 140
rect -3915 50 -3875 60
rect -3825 140 -3785 150
rect -3825 60 -3815 140
rect -3795 60 -3785 140
rect -3825 50 -3785 60
rect -3735 140 -3695 150
rect -3735 60 -3725 140
rect -3705 60 -3695 140
rect -3735 50 -3695 60
rect -3645 140 -3605 150
rect -3645 60 -3635 140
rect -3615 60 -3605 140
rect -3645 50 -3605 60
rect -3555 140 -3515 150
rect -3555 60 -3545 140
rect -3525 60 -3515 140
rect -3555 50 -3515 60
rect -3465 140 -3425 150
rect -3465 60 -3455 140
rect -3435 60 -3425 140
rect -3465 50 -3425 60
rect -3375 140 -3335 150
rect -3375 60 -3365 140
rect -3345 60 -3335 140
rect -3375 50 -3335 60
rect -3285 140 -3245 150
rect -3285 60 -3275 140
rect -3255 60 -3245 140
rect -3285 50 -3245 60
rect -3195 140 -3155 150
rect -3195 60 -3185 140
rect -3165 60 -3155 140
rect -3195 50 -3155 60
rect -3105 140 -3065 150
rect -3105 60 -3095 140
rect -3075 60 -3065 140
rect -3105 50 -3065 60
rect -3015 140 -2975 150
rect -3015 60 -3005 140
rect -2985 60 -2975 140
rect -3015 50 -2975 60
rect -2925 140 -2885 150
rect -2925 60 -2915 140
rect -2895 60 -2885 140
rect -2925 50 -2885 60
rect -2835 140 -2795 150
rect -2835 60 -2825 140
rect -2805 60 -2795 140
rect -2835 50 -2795 60
rect -2745 140 -2705 150
rect -2745 60 -2735 140
rect -2715 60 -2705 140
rect -2745 50 -2705 60
rect -2655 140 -2615 150
rect -2655 60 -2645 140
rect -2625 60 -2615 140
rect -2655 50 -2615 60
rect -2565 140 -2525 150
rect -2565 60 -2555 140
rect -2535 60 -2525 140
rect -2565 50 -2525 60
rect -2475 140 -2435 150
rect -2475 60 -2465 140
rect -2445 60 -2435 140
rect -2475 50 -2435 60
rect -2385 140 -2345 150
rect -2385 60 -2375 140
rect -2355 60 -2345 140
rect -2385 50 -2345 60
rect -2295 140 -2255 150
rect -2295 60 -2285 140
rect -2265 60 -2255 140
rect -2295 50 -2255 60
rect -2205 140 -2165 150
rect -2205 60 -2195 140
rect -2175 60 -2165 140
rect -2205 50 -2165 60
rect -2115 140 -2075 150
rect -2115 60 -2105 140
rect -2085 60 -2075 140
rect -2115 50 -2075 60
rect -2025 140 -1985 150
rect -2025 60 -2015 140
rect -1995 60 -1985 140
rect -2025 50 -1985 60
rect -1935 140 -1895 150
rect -1935 60 -1925 140
rect -1905 60 -1895 140
rect -1935 50 -1895 60
rect -1845 140 -1805 150
rect -1845 60 -1835 140
rect -1815 60 -1805 140
rect -1845 50 -1805 60
rect -1755 140 -1715 150
rect -1755 60 -1745 140
rect -1725 60 -1715 140
rect -1755 50 -1715 60
rect -1665 140 -1625 150
rect -1665 60 -1655 140
rect -1635 60 -1625 140
rect -1665 50 -1625 60
rect -1575 140 -1535 150
rect -1575 60 -1565 140
rect -1545 60 -1535 140
rect -1575 50 -1535 60
rect -1485 140 -1445 150
rect -1485 60 -1475 140
rect -1455 60 -1445 140
rect -1485 50 -1445 60
rect -1395 140 -1355 150
rect -1395 60 -1385 140
rect -1365 60 -1355 140
rect -1395 50 -1355 60
rect -1305 140 -1265 150
rect -1305 60 -1295 140
rect -1275 60 -1265 140
rect -1305 50 -1265 60
rect -1215 140 -1175 150
rect -1215 60 -1205 140
rect -1185 60 -1175 140
rect -1215 50 -1175 60
rect -1125 140 -1085 150
rect -1125 60 -1115 140
rect -1095 60 -1085 140
rect -1125 50 -1085 60
rect -1035 140 -995 150
rect -1035 60 -1025 140
rect -1005 60 -995 140
rect -1035 50 -995 60
rect -945 140 -905 150
rect -945 60 -935 140
rect -915 60 -905 140
rect -945 50 -905 60
rect -855 140 -815 150
rect -855 60 -845 140
rect -825 60 -815 140
rect -855 50 -815 60
rect -765 140 -725 150
rect -765 60 -755 140
rect -735 60 -725 140
rect -765 50 -725 60
rect -675 140 -635 150
rect -675 60 -665 140
rect -645 60 -635 140
rect -675 50 -635 60
rect -585 140 -545 150
rect -585 60 -575 140
rect -555 60 -545 140
rect -585 50 -545 60
rect -495 140 -455 150
rect -495 60 -485 140
rect -465 60 -455 140
rect -495 50 -455 60
rect -405 140 -365 150
rect -405 60 -395 140
rect -375 60 -365 140
rect -405 50 -365 60
rect -315 140 -275 150
rect -315 60 -305 140
rect -285 60 -275 140
rect -315 50 -275 60
rect -225 140 -185 150
rect -225 60 -215 140
rect -195 60 -185 140
rect -225 50 -185 60
rect -135 140 -95 150
rect -135 60 -125 140
rect -105 60 -95 140
rect -135 50 -95 60
rect -45 140 -5 150
rect -45 60 -35 140
rect -15 60 -5 140
rect -45 50 -5 60
<< mvpdiff >>
rect -11565 1155 -11525 1165
rect -11565 1075 -11555 1155
rect -11535 1075 -11525 1155
rect -11565 1065 -11525 1075
rect -11475 1155 -11435 1165
rect -11475 1075 -11465 1155
rect -11445 1075 -11435 1155
rect -11475 1065 -11435 1075
rect -11385 1155 -11345 1165
rect -11385 1075 -11375 1155
rect -11355 1075 -11345 1155
rect -11385 1065 -11345 1075
rect -11295 1155 -11255 1165
rect -11295 1075 -11285 1155
rect -11265 1075 -11255 1155
rect -11295 1065 -11255 1075
rect -11205 1155 -11165 1165
rect -11205 1075 -11195 1155
rect -11175 1075 -11165 1155
rect -11205 1065 -11165 1075
rect -11115 1155 -11075 1165
rect -11115 1075 -11105 1155
rect -11085 1075 -11075 1155
rect -11115 1065 -11075 1075
rect -11025 1155 -10985 1165
rect -11025 1075 -11015 1155
rect -10995 1075 -10985 1155
rect -11025 1065 -10985 1075
rect -10935 1155 -10895 1165
rect -10935 1075 -10925 1155
rect -10905 1075 -10895 1155
rect -10935 1065 -10895 1075
rect -10845 1155 -10805 1165
rect -10845 1075 -10835 1155
rect -10815 1075 -10805 1155
rect -10845 1065 -10805 1075
rect -10755 1155 -10715 1165
rect -10755 1075 -10745 1155
rect -10725 1075 -10715 1155
rect -10755 1065 -10715 1075
rect -10665 1155 -10625 1165
rect -10665 1075 -10655 1155
rect -10635 1075 -10625 1155
rect -10665 1065 -10625 1075
rect -10575 1155 -10535 1165
rect -10575 1075 -10565 1155
rect -10545 1075 -10535 1155
rect -10575 1065 -10535 1075
rect -10485 1155 -10445 1165
rect -10485 1075 -10475 1155
rect -10455 1075 -10445 1155
rect -10485 1065 -10445 1075
rect -10395 1155 -10355 1165
rect -10395 1075 -10385 1155
rect -10365 1075 -10355 1155
rect -10395 1065 -10355 1075
rect -10305 1155 -10265 1165
rect -10305 1075 -10295 1155
rect -10275 1075 -10265 1155
rect -10305 1065 -10265 1075
rect -10215 1155 -10175 1165
rect -10215 1075 -10205 1155
rect -10185 1075 -10175 1155
rect -10215 1065 -10175 1075
rect -10125 1155 -10085 1165
rect -10125 1075 -10115 1155
rect -10095 1075 -10085 1155
rect -10125 1065 -10085 1075
rect -10035 1155 -9995 1165
rect -10035 1075 -10025 1155
rect -10005 1075 -9995 1155
rect -10035 1065 -9995 1075
rect -9945 1155 -9905 1165
rect -9945 1075 -9935 1155
rect -9915 1075 -9905 1155
rect -9945 1065 -9905 1075
rect -9855 1155 -9815 1165
rect -9855 1075 -9845 1155
rect -9825 1075 -9815 1155
rect -9855 1065 -9815 1075
rect -9765 1155 -9725 1165
rect -9765 1075 -9755 1155
rect -9735 1075 -9725 1155
rect -9765 1065 -9725 1075
rect -9675 1155 -9635 1165
rect -9675 1075 -9665 1155
rect -9645 1075 -9635 1155
rect -9675 1065 -9635 1075
rect -9585 1155 -9545 1165
rect -9585 1075 -9575 1155
rect -9555 1075 -9545 1155
rect -9585 1065 -9545 1075
rect -9495 1155 -9455 1165
rect -9495 1075 -9485 1155
rect -9465 1075 -9455 1155
rect -9495 1065 -9455 1075
rect -9405 1155 -9365 1165
rect -9405 1075 -9395 1155
rect -9375 1075 -9365 1155
rect -9405 1065 -9365 1075
rect -9315 1155 -9275 1165
rect -9315 1075 -9305 1155
rect -9285 1075 -9275 1155
rect -9315 1065 -9275 1075
rect -9225 1155 -9185 1165
rect -9225 1075 -9215 1155
rect -9195 1075 -9185 1155
rect -9225 1065 -9185 1075
rect -9135 1155 -9095 1165
rect -9135 1075 -9125 1155
rect -9105 1075 -9095 1155
rect -9135 1065 -9095 1075
rect -9045 1155 -9005 1165
rect -9045 1075 -9035 1155
rect -9015 1075 -9005 1155
rect -9045 1065 -9005 1075
rect -8955 1155 -8915 1165
rect -8955 1075 -8945 1155
rect -8925 1075 -8915 1155
rect -8955 1065 -8915 1075
rect -8865 1155 -8825 1165
rect -8865 1075 -8855 1155
rect -8835 1075 -8825 1155
rect -8865 1065 -8825 1075
rect -8775 1155 -8735 1165
rect -8775 1075 -8765 1155
rect -8745 1075 -8735 1155
rect -8775 1065 -8735 1075
rect -8685 1155 -8645 1165
rect -8685 1075 -8675 1155
rect -8655 1075 -8645 1155
rect -8685 1065 -8645 1075
rect -8595 1155 -8555 1165
rect -8595 1075 -8585 1155
rect -8565 1075 -8555 1155
rect -8595 1065 -8555 1075
rect -8505 1155 -8465 1165
rect -8505 1075 -8495 1155
rect -8475 1075 -8465 1155
rect -8505 1065 -8465 1075
rect -8415 1155 -8375 1165
rect -8415 1075 -8405 1155
rect -8385 1075 -8375 1155
rect -8415 1065 -8375 1075
rect -8325 1155 -8285 1165
rect -8325 1075 -8315 1155
rect -8295 1075 -8285 1155
rect -8325 1065 -8285 1075
rect -8235 1155 -8195 1165
rect -8235 1075 -8225 1155
rect -8205 1075 -8195 1155
rect -8235 1065 -8195 1075
rect -8145 1155 -8105 1165
rect -8145 1075 -8135 1155
rect -8115 1075 -8105 1155
rect -8145 1065 -8105 1075
rect -8055 1155 -8015 1165
rect -8055 1075 -8045 1155
rect -8025 1075 -8015 1155
rect -8055 1065 -8015 1075
rect -7965 1155 -7925 1165
rect -7965 1075 -7955 1155
rect -7935 1075 -7925 1155
rect -7965 1065 -7925 1075
rect -7875 1155 -7835 1165
rect -7875 1075 -7865 1155
rect -7845 1075 -7835 1155
rect -7875 1065 -7835 1075
rect -7785 1155 -7745 1165
rect -7785 1075 -7775 1155
rect -7755 1075 -7745 1155
rect -7785 1065 -7745 1075
rect -7695 1155 -7655 1165
rect -7695 1075 -7685 1155
rect -7665 1075 -7655 1155
rect -7695 1065 -7655 1075
rect -7605 1155 -7565 1165
rect -7605 1075 -7595 1155
rect -7575 1075 -7565 1155
rect -7605 1065 -7565 1075
rect -7515 1155 -7475 1165
rect -7515 1075 -7505 1155
rect -7485 1075 -7475 1155
rect -7515 1065 -7475 1075
rect -7425 1155 -7385 1165
rect -7425 1075 -7415 1155
rect -7395 1075 -7385 1155
rect -7425 1065 -7385 1075
rect -7335 1155 -7295 1165
rect -7335 1075 -7325 1155
rect -7305 1075 -7295 1155
rect -7335 1065 -7295 1075
rect -7245 1155 -7205 1165
rect -7245 1075 -7235 1155
rect -7215 1075 -7205 1155
rect -7245 1065 -7205 1075
rect -7155 1155 -7115 1165
rect -7155 1075 -7145 1155
rect -7125 1075 -7115 1155
rect -7155 1065 -7115 1075
rect -7065 1155 -7025 1165
rect -7065 1075 -7055 1155
rect -7035 1075 -7025 1155
rect -7065 1065 -7025 1075
rect -6975 1155 -6935 1165
rect -6975 1075 -6965 1155
rect -6945 1075 -6935 1155
rect -6975 1065 -6935 1075
rect -6885 1155 -6845 1165
rect -6885 1075 -6875 1155
rect -6855 1075 -6845 1155
rect -6885 1065 -6845 1075
rect -6795 1155 -6755 1165
rect -6795 1075 -6785 1155
rect -6765 1075 -6755 1155
rect -6795 1065 -6755 1075
rect -6705 1155 -6665 1165
rect -6705 1075 -6695 1155
rect -6675 1075 -6665 1155
rect -6705 1065 -6665 1075
rect -6615 1155 -6575 1165
rect -6615 1075 -6605 1155
rect -6585 1075 -6575 1155
rect -6615 1065 -6575 1075
rect -6525 1155 -6485 1165
rect -6525 1075 -6515 1155
rect -6495 1075 -6485 1155
rect -6525 1065 -6485 1075
rect -6435 1155 -6395 1165
rect -6435 1075 -6425 1155
rect -6405 1075 -6395 1155
rect -6435 1065 -6395 1075
rect -6345 1155 -6305 1165
rect -6345 1075 -6335 1155
rect -6315 1075 -6305 1155
rect -6345 1065 -6305 1075
rect -6255 1155 -6215 1165
rect -6255 1075 -6245 1155
rect -6225 1075 -6215 1155
rect -6255 1065 -6215 1075
rect -6165 1155 -6125 1165
rect -6165 1075 -6155 1155
rect -6135 1075 -6125 1155
rect -6165 1065 -6125 1075
rect -6075 1155 -6035 1165
rect -6075 1075 -6065 1155
rect -6045 1075 -6035 1155
rect -6075 1065 -6035 1075
rect -5985 1155 -5945 1165
rect -5985 1075 -5975 1155
rect -5955 1075 -5945 1155
rect -5985 1065 -5945 1075
rect -5895 1155 -5855 1165
rect -5895 1075 -5885 1155
rect -5865 1075 -5855 1155
rect -5895 1065 -5855 1075
rect -5805 1155 -5765 1165
rect -5805 1075 -5795 1155
rect -5775 1075 -5765 1155
rect -5805 1065 -5765 1075
rect -5715 1155 -5675 1165
rect -5715 1075 -5705 1155
rect -5685 1075 -5675 1155
rect -5715 1065 -5675 1075
rect -5625 1155 -5585 1165
rect -5625 1075 -5615 1155
rect -5595 1075 -5585 1155
rect -5625 1065 -5585 1075
rect -5535 1155 -5495 1165
rect -5535 1075 -5525 1155
rect -5505 1075 -5495 1155
rect -5535 1065 -5495 1075
rect -5445 1155 -5405 1165
rect -5445 1075 -5435 1155
rect -5415 1075 -5405 1155
rect -5445 1065 -5405 1075
rect -5355 1155 -5315 1165
rect -5355 1075 -5345 1155
rect -5325 1075 -5315 1155
rect -5355 1065 -5315 1075
rect -5265 1155 -5225 1165
rect -5265 1075 -5255 1155
rect -5235 1075 -5225 1155
rect -5265 1065 -5225 1075
rect -5175 1155 -5135 1165
rect -5175 1075 -5165 1155
rect -5145 1075 -5135 1155
rect -5175 1065 -5135 1075
rect -5085 1155 -5045 1165
rect -5085 1075 -5075 1155
rect -5055 1075 -5045 1155
rect -5085 1065 -5045 1075
rect -4995 1155 -4955 1165
rect -4995 1075 -4985 1155
rect -4965 1075 -4955 1155
rect -4995 1065 -4955 1075
rect -4905 1155 -4865 1165
rect -4905 1075 -4895 1155
rect -4875 1075 -4865 1155
rect -4905 1065 -4865 1075
rect -4815 1155 -4775 1165
rect -4815 1075 -4805 1155
rect -4785 1075 -4775 1155
rect -4815 1065 -4775 1075
rect -4725 1155 -4685 1165
rect -4725 1075 -4715 1155
rect -4695 1075 -4685 1155
rect -4725 1065 -4685 1075
rect -4635 1155 -4595 1165
rect -4635 1075 -4625 1155
rect -4605 1075 -4595 1155
rect -4635 1065 -4595 1075
rect -4545 1155 -4505 1165
rect -4545 1075 -4535 1155
rect -4515 1075 -4505 1155
rect -4545 1065 -4505 1075
rect -4455 1155 -4415 1165
rect -4455 1075 -4445 1155
rect -4425 1075 -4415 1155
rect -4455 1065 -4415 1075
rect -4365 1155 -4325 1165
rect -4365 1075 -4355 1155
rect -4335 1075 -4325 1155
rect -4365 1065 -4325 1075
rect -4275 1155 -4235 1165
rect -4275 1075 -4265 1155
rect -4245 1075 -4235 1155
rect -4275 1065 -4235 1075
rect -4185 1155 -4145 1165
rect -4185 1075 -4175 1155
rect -4155 1075 -4145 1155
rect -4185 1065 -4145 1075
rect -4095 1155 -4055 1165
rect -4095 1075 -4085 1155
rect -4065 1075 -4055 1155
rect -4095 1065 -4055 1075
rect -4005 1155 -3965 1165
rect -4005 1075 -3995 1155
rect -3975 1075 -3965 1155
rect -4005 1065 -3965 1075
rect -3915 1155 -3875 1165
rect -3915 1075 -3905 1155
rect -3885 1075 -3875 1155
rect -3915 1065 -3875 1075
rect -3825 1155 -3785 1165
rect -3825 1075 -3815 1155
rect -3795 1075 -3785 1155
rect -3825 1065 -3785 1075
rect -3735 1155 -3695 1165
rect -3735 1075 -3725 1155
rect -3705 1075 -3695 1155
rect -3735 1065 -3695 1075
rect -3645 1155 -3605 1165
rect -3645 1075 -3635 1155
rect -3615 1075 -3605 1155
rect -3645 1065 -3605 1075
rect -3555 1155 -3515 1165
rect -3555 1075 -3545 1155
rect -3525 1075 -3515 1155
rect -3555 1065 -3515 1075
rect -3465 1155 -3425 1165
rect -3465 1075 -3455 1155
rect -3435 1075 -3425 1155
rect -3465 1065 -3425 1075
rect -3375 1155 -3335 1165
rect -3375 1075 -3365 1155
rect -3345 1075 -3335 1155
rect -3375 1065 -3335 1075
rect -3285 1155 -3245 1165
rect -3285 1075 -3275 1155
rect -3255 1075 -3245 1155
rect -3285 1065 -3245 1075
rect -3195 1155 -3155 1165
rect -3195 1075 -3185 1155
rect -3165 1075 -3155 1155
rect -3195 1065 -3155 1075
rect -3105 1155 -3065 1165
rect -3105 1075 -3095 1155
rect -3075 1075 -3065 1155
rect -3105 1065 -3065 1075
rect -3015 1155 -2975 1165
rect -3015 1075 -3005 1155
rect -2985 1075 -2975 1155
rect -3015 1065 -2975 1075
rect -2925 1155 -2885 1165
rect -2925 1075 -2915 1155
rect -2895 1075 -2885 1155
rect -2925 1065 -2885 1075
rect -2835 1155 -2795 1165
rect -2835 1075 -2825 1155
rect -2805 1075 -2795 1155
rect -2835 1065 -2795 1075
rect -2745 1155 -2705 1165
rect -2745 1075 -2735 1155
rect -2715 1075 -2705 1155
rect -2745 1065 -2705 1075
rect -2655 1155 -2615 1165
rect -2655 1075 -2645 1155
rect -2625 1075 -2615 1155
rect -2655 1065 -2615 1075
rect -2565 1155 -2525 1165
rect -2565 1075 -2555 1155
rect -2535 1075 -2525 1155
rect -2565 1065 -2525 1075
rect -2475 1155 -2435 1165
rect -2475 1075 -2465 1155
rect -2445 1075 -2435 1155
rect -2475 1065 -2435 1075
rect -2385 1155 -2345 1165
rect -2385 1075 -2375 1155
rect -2355 1075 -2345 1155
rect -2385 1065 -2345 1075
rect -2295 1155 -2255 1165
rect -2295 1075 -2285 1155
rect -2265 1075 -2255 1155
rect -2295 1065 -2255 1075
rect -2205 1155 -2165 1165
rect -2205 1075 -2195 1155
rect -2175 1075 -2165 1155
rect -2205 1065 -2165 1075
rect -2115 1155 -2075 1165
rect -2115 1075 -2105 1155
rect -2085 1075 -2075 1155
rect -2115 1065 -2075 1075
rect -2025 1155 -1985 1165
rect -2025 1075 -2015 1155
rect -1995 1075 -1985 1155
rect -2025 1065 -1985 1075
rect -1935 1155 -1895 1165
rect -1935 1075 -1925 1155
rect -1905 1075 -1895 1155
rect -1935 1065 -1895 1075
rect -1845 1155 -1805 1165
rect -1845 1075 -1835 1155
rect -1815 1075 -1805 1155
rect -1845 1065 -1805 1075
rect -1755 1155 -1715 1165
rect -1755 1075 -1745 1155
rect -1725 1075 -1715 1155
rect -1755 1065 -1715 1075
rect -1665 1155 -1625 1165
rect -1665 1075 -1655 1155
rect -1635 1075 -1625 1155
rect -1665 1065 -1625 1075
rect -1575 1155 -1535 1165
rect -1575 1075 -1565 1155
rect -1545 1075 -1535 1155
rect -1575 1065 -1535 1075
rect -1485 1155 -1445 1165
rect -1485 1075 -1475 1155
rect -1455 1075 -1445 1155
rect -1485 1065 -1445 1075
rect -1395 1155 -1355 1165
rect -1395 1075 -1385 1155
rect -1365 1075 -1355 1155
rect -1395 1065 -1355 1075
rect -1305 1155 -1265 1165
rect -1305 1075 -1295 1155
rect -1275 1075 -1265 1155
rect -1305 1065 -1265 1075
rect -1215 1155 -1175 1165
rect -1215 1075 -1205 1155
rect -1185 1075 -1175 1155
rect -1215 1065 -1175 1075
rect -1125 1155 -1085 1165
rect -1125 1075 -1115 1155
rect -1095 1075 -1085 1155
rect -1125 1065 -1085 1075
rect -1035 1155 -995 1165
rect -1035 1075 -1025 1155
rect -1005 1075 -995 1155
rect -1035 1065 -995 1075
rect -945 1155 -905 1165
rect -945 1075 -935 1155
rect -915 1075 -905 1155
rect -945 1065 -905 1075
rect -855 1155 -815 1165
rect -855 1075 -845 1155
rect -825 1075 -815 1155
rect -855 1065 -815 1075
rect -765 1155 -725 1165
rect -765 1075 -755 1155
rect -735 1075 -725 1155
rect -765 1065 -725 1075
rect -675 1155 -635 1165
rect -675 1075 -665 1155
rect -645 1075 -635 1155
rect -675 1065 -635 1075
rect -585 1155 -545 1165
rect -585 1075 -575 1155
rect -555 1075 -545 1155
rect -585 1065 -545 1075
rect -495 1155 -455 1165
rect -495 1075 -485 1155
rect -465 1075 -455 1155
rect -495 1065 -455 1075
rect -405 1155 -365 1165
rect -405 1075 -395 1155
rect -375 1075 -365 1155
rect -405 1065 -365 1075
rect -315 1155 -275 1165
rect -315 1075 -305 1155
rect -285 1075 -275 1155
rect -315 1065 -275 1075
rect -225 1155 -185 1165
rect -225 1075 -215 1155
rect -195 1075 -185 1155
rect -225 1065 -185 1075
rect -135 1155 -95 1165
rect -135 1075 -125 1155
rect -105 1075 -95 1155
rect -135 1065 -95 1075
rect -45 1155 -5 1165
rect -45 1075 -35 1155
rect -15 1075 -5 1155
rect -45 1065 -5 1075
rect -11565 920 -11525 930
rect -11565 840 -11555 920
rect -11535 840 -11525 920
rect -11565 830 -11525 840
rect -11475 920 -11435 930
rect -11475 840 -11465 920
rect -11445 840 -11435 920
rect -11475 830 -11435 840
rect -11385 920 -11345 930
rect -11385 840 -11375 920
rect -11355 840 -11345 920
rect -11385 830 -11345 840
rect -11295 920 -11255 930
rect -11295 840 -11285 920
rect -11265 840 -11255 920
rect -11295 830 -11255 840
rect -11205 920 -11165 930
rect -11205 840 -11195 920
rect -11175 840 -11165 920
rect -11205 830 -11165 840
rect -11115 920 -11075 930
rect -11115 840 -11105 920
rect -11085 840 -11075 920
rect -11115 830 -11075 840
rect -11025 920 -10985 930
rect -11025 840 -11015 920
rect -10995 840 -10985 920
rect -11025 830 -10985 840
rect -10935 920 -10895 930
rect -10935 840 -10925 920
rect -10905 840 -10895 920
rect -10935 830 -10895 840
rect -10845 920 -10805 930
rect -10845 840 -10835 920
rect -10815 840 -10805 920
rect -10845 830 -10805 840
rect -10755 920 -10715 930
rect -10755 840 -10745 920
rect -10725 840 -10715 920
rect -10755 830 -10715 840
rect -10665 920 -10625 930
rect -10665 840 -10655 920
rect -10635 840 -10625 920
rect -10665 830 -10625 840
rect -10575 920 -10535 930
rect -10575 840 -10565 920
rect -10545 840 -10535 920
rect -10575 830 -10535 840
rect -10485 920 -10445 930
rect -10485 840 -10475 920
rect -10455 840 -10445 920
rect -10485 830 -10445 840
rect -10395 920 -10355 930
rect -10395 840 -10385 920
rect -10365 840 -10355 920
rect -10395 830 -10355 840
rect -10305 920 -10265 930
rect -10305 840 -10295 920
rect -10275 840 -10265 920
rect -10305 830 -10265 840
rect -10215 920 -10175 930
rect -10215 840 -10205 920
rect -10185 840 -10175 920
rect -10215 830 -10175 840
rect -10125 920 -10085 930
rect -10125 840 -10115 920
rect -10095 840 -10085 920
rect -10125 830 -10085 840
rect -10035 920 -9995 930
rect -10035 840 -10025 920
rect -10005 840 -9995 920
rect -10035 830 -9995 840
rect -9945 920 -9905 930
rect -9945 840 -9935 920
rect -9915 840 -9905 920
rect -9945 830 -9905 840
rect -9855 920 -9815 930
rect -9855 840 -9845 920
rect -9825 840 -9815 920
rect -9855 830 -9815 840
rect -9765 920 -9725 930
rect -9765 840 -9755 920
rect -9735 840 -9725 920
rect -9765 830 -9725 840
rect -9675 920 -9635 930
rect -9675 840 -9665 920
rect -9645 840 -9635 920
rect -9675 830 -9635 840
rect -9585 920 -9545 930
rect -9585 840 -9575 920
rect -9555 840 -9545 920
rect -9585 830 -9545 840
rect -9495 920 -9455 930
rect -9495 840 -9485 920
rect -9465 840 -9455 920
rect -9495 830 -9455 840
rect -9405 920 -9365 930
rect -9405 840 -9395 920
rect -9375 840 -9365 920
rect -9405 830 -9365 840
rect -9315 920 -9275 930
rect -9315 840 -9305 920
rect -9285 840 -9275 920
rect -9315 830 -9275 840
rect -9225 920 -9185 930
rect -9225 840 -9215 920
rect -9195 840 -9185 920
rect -9225 830 -9185 840
rect -9135 920 -9095 930
rect -9135 840 -9125 920
rect -9105 840 -9095 920
rect -9135 830 -9095 840
rect -9045 920 -9005 930
rect -9045 840 -9035 920
rect -9015 840 -9005 920
rect -9045 830 -9005 840
rect -8955 920 -8915 930
rect -8955 840 -8945 920
rect -8925 840 -8915 920
rect -8955 830 -8915 840
rect -8865 920 -8825 930
rect -8865 840 -8855 920
rect -8835 840 -8825 920
rect -8865 830 -8825 840
rect -8775 920 -8735 930
rect -8775 840 -8765 920
rect -8745 840 -8735 920
rect -8775 830 -8735 840
rect -8685 920 -8645 930
rect -8685 840 -8675 920
rect -8655 840 -8645 920
rect -8685 830 -8645 840
rect -8595 920 -8555 930
rect -8595 840 -8585 920
rect -8565 840 -8555 920
rect -8595 830 -8555 840
rect -8505 920 -8465 930
rect -8505 840 -8495 920
rect -8475 840 -8465 920
rect -8505 830 -8465 840
rect -8415 920 -8375 930
rect -8415 840 -8405 920
rect -8385 840 -8375 920
rect -8415 830 -8375 840
rect -8325 920 -8285 930
rect -8325 840 -8315 920
rect -8295 840 -8285 920
rect -8325 830 -8285 840
rect -8235 920 -8195 930
rect -8235 840 -8225 920
rect -8205 840 -8195 920
rect -8235 830 -8195 840
rect -8145 920 -8105 930
rect -8145 840 -8135 920
rect -8115 840 -8105 920
rect -8145 830 -8105 840
rect -8055 920 -8015 930
rect -8055 840 -8045 920
rect -8025 840 -8015 920
rect -8055 830 -8015 840
rect -7965 920 -7925 930
rect -7965 840 -7955 920
rect -7935 840 -7925 920
rect -7965 830 -7925 840
rect -7875 920 -7835 930
rect -7875 840 -7865 920
rect -7845 840 -7835 920
rect -7875 830 -7835 840
rect -7785 920 -7745 930
rect -7785 840 -7775 920
rect -7755 840 -7745 920
rect -7785 830 -7745 840
rect -7695 920 -7655 930
rect -7695 840 -7685 920
rect -7665 840 -7655 920
rect -7695 830 -7655 840
rect -7605 920 -7565 930
rect -7605 840 -7595 920
rect -7575 840 -7565 920
rect -7605 830 -7565 840
rect -7515 920 -7475 930
rect -7515 840 -7505 920
rect -7485 840 -7475 920
rect -7515 830 -7475 840
rect -7425 920 -7385 930
rect -7425 840 -7415 920
rect -7395 840 -7385 920
rect -7425 830 -7385 840
rect -7335 920 -7295 930
rect -7335 840 -7325 920
rect -7305 840 -7295 920
rect -7335 830 -7295 840
rect -7245 920 -7205 930
rect -7245 840 -7235 920
rect -7215 840 -7205 920
rect -7245 830 -7205 840
rect -7155 920 -7115 930
rect -7155 840 -7145 920
rect -7125 840 -7115 920
rect -7155 830 -7115 840
rect -7065 920 -7025 930
rect -7065 840 -7055 920
rect -7035 840 -7025 920
rect -7065 830 -7025 840
rect -6975 920 -6935 930
rect -6975 840 -6965 920
rect -6945 840 -6935 920
rect -6975 830 -6935 840
rect -6885 920 -6845 930
rect -6885 840 -6875 920
rect -6855 840 -6845 920
rect -6885 830 -6845 840
rect -6795 920 -6755 930
rect -6795 840 -6785 920
rect -6765 840 -6755 920
rect -6795 830 -6755 840
rect -6705 920 -6665 930
rect -6705 840 -6695 920
rect -6675 840 -6665 920
rect -6705 830 -6665 840
rect -6615 920 -6575 930
rect -6615 840 -6605 920
rect -6585 840 -6575 920
rect -6615 830 -6575 840
rect -6525 920 -6485 930
rect -6525 840 -6515 920
rect -6495 840 -6485 920
rect -6525 830 -6485 840
rect -6435 920 -6395 930
rect -6435 840 -6425 920
rect -6405 840 -6395 920
rect -6435 830 -6395 840
rect -6345 920 -6305 930
rect -6345 840 -6335 920
rect -6315 840 -6305 920
rect -6345 830 -6305 840
rect -6255 920 -6215 930
rect -6255 840 -6245 920
rect -6225 840 -6215 920
rect -6255 830 -6215 840
rect -6165 920 -6125 930
rect -6165 840 -6155 920
rect -6135 840 -6125 920
rect -6165 830 -6125 840
rect -6075 920 -6035 930
rect -6075 840 -6065 920
rect -6045 840 -6035 920
rect -6075 830 -6035 840
rect -5985 920 -5945 930
rect -5985 840 -5975 920
rect -5955 840 -5945 920
rect -5985 830 -5945 840
rect -5895 920 -5855 930
rect -5895 840 -5885 920
rect -5865 840 -5855 920
rect -5895 830 -5855 840
rect -5805 920 -5765 930
rect -5805 840 -5795 920
rect -5775 840 -5765 920
rect -5805 830 -5765 840
rect -5715 920 -5675 930
rect -5715 840 -5705 920
rect -5685 840 -5675 920
rect -5715 830 -5675 840
rect -5625 920 -5585 930
rect -5625 840 -5615 920
rect -5595 840 -5585 920
rect -5625 830 -5585 840
rect -5535 920 -5495 930
rect -5535 840 -5525 920
rect -5505 840 -5495 920
rect -5535 830 -5495 840
rect -5445 920 -5405 930
rect -5445 840 -5435 920
rect -5415 840 -5405 920
rect -5445 830 -5405 840
rect -5355 920 -5315 930
rect -5355 840 -5345 920
rect -5325 840 -5315 920
rect -5355 830 -5315 840
rect -5265 920 -5225 930
rect -5265 840 -5255 920
rect -5235 840 -5225 920
rect -5265 830 -5225 840
rect -5175 920 -5135 930
rect -5175 840 -5165 920
rect -5145 840 -5135 920
rect -5175 830 -5135 840
rect -5085 920 -5045 930
rect -5085 840 -5075 920
rect -5055 840 -5045 920
rect -5085 830 -5045 840
rect -4995 920 -4955 930
rect -4995 840 -4985 920
rect -4965 840 -4955 920
rect -4995 830 -4955 840
rect -4905 920 -4865 930
rect -4905 840 -4895 920
rect -4875 840 -4865 920
rect -4905 830 -4865 840
rect -4815 920 -4775 930
rect -4815 840 -4805 920
rect -4785 840 -4775 920
rect -4815 830 -4775 840
rect -4725 920 -4685 930
rect -4725 840 -4715 920
rect -4695 840 -4685 920
rect -4725 830 -4685 840
rect -4635 920 -4595 930
rect -4635 840 -4625 920
rect -4605 840 -4595 920
rect -4635 830 -4595 840
rect -4545 920 -4505 930
rect -4545 840 -4535 920
rect -4515 840 -4505 920
rect -4545 830 -4505 840
rect -4455 920 -4415 930
rect -4455 840 -4445 920
rect -4425 840 -4415 920
rect -4455 830 -4415 840
rect -4365 920 -4325 930
rect -4365 840 -4355 920
rect -4335 840 -4325 920
rect -4365 830 -4325 840
rect -4275 920 -4235 930
rect -4275 840 -4265 920
rect -4245 840 -4235 920
rect -4275 830 -4235 840
rect -4185 920 -4145 930
rect -4185 840 -4175 920
rect -4155 840 -4145 920
rect -4185 830 -4145 840
rect -4095 920 -4055 930
rect -4095 840 -4085 920
rect -4065 840 -4055 920
rect -4095 830 -4055 840
rect -4005 920 -3965 930
rect -4005 840 -3995 920
rect -3975 840 -3965 920
rect -4005 830 -3965 840
rect -3915 920 -3875 930
rect -3915 840 -3905 920
rect -3885 840 -3875 920
rect -3915 830 -3875 840
rect -3825 920 -3785 930
rect -3825 840 -3815 920
rect -3795 840 -3785 920
rect -3825 830 -3785 840
rect -3735 920 -3695 930
rect -3735 840 -3725 920
rect -3705 840 -3695 920
rect -3735 830 -3695 840
rect -3645 920 -3605 930
rect -3645 840 -3635 920
rect -3615 840 -3605 920
rect -3645 830 -3605 840
rect -3555 920 -3515 930
rect -3555 840 -3545 920
rect -3525 840 -3515 920
rect -3555 830 -3515 840
rect -3465 920 -3425 930
rect -3465 840 -3455 920
rect -3435 840 -3425 920
rect -3465 830 -3425 840
rect -3375 920 -3335 930
rect -3375 840 -3365 920
rect -3345 840 -3335 920
rect -3375 830 -3335 840
rect -3285 920 -3245 930
rect -3285 840 -3275 920
rect -3255 840 -3245 920
rect -3285 830 -3245 840
rect -3195 920 -3155 930
rect -3195 840 -3185 920
rect -3165 840 -3155 920
rect -3195 830 -3155 840
rect -3105 920 -3065 930
rect -3105 840 -3095 920
rect -3075 840 -3065 920
rect -3105 830 -3065 840
rect -3015 920 -2975 930
rect -3015 840 -3005 920
rect -2985 840 -2975 920
rect -3015 830 -2975 840
rect -2925 920 -2885 930
rect -2925 840 -2915 920
rect -2895 840 -2885 920
rect -2925 830 -2885 840
rect -2835 920 -2795 930
rect -2835 840 -2825 920
rect -2805 840 -2795 920
rect -2835 830 -2795 840
rect -2745 920 -2705 930
rect -2745 840 -2735 920
rect -2715 840 -2705 920
rect -2745 830 -2705 840
rect -2655 920 -2615 930
rect -2655 840 -2645 920
rect -2625 840 -2615 920
rect -2655 830 -2615 840
rect -2565 920 -2525 930
rect -2565 840 -2555 920
rect -2535 840 -2525 920
rect -2565 830 -2525 840
rect -2475 920 -2435 930
rect -2475 840 -2465 920
rect -2445 840 -2435 920
rect -2475 830 -2435 840
rect -2385 920 -2345 930
rect -2385 840 -2375 920
rect -2355 840 -2345 920
rect -2385 830 -2345 840
rect -2295 920 -2255 930
rect -2295 840 -2285 920
rect -2265 840 -2255 920
rect -2295 830 -2255 840
rect -2205 920 -2165 930
rect -2205 840 -2195 920
rect -2175 840 -2165 920
rect -2205 830 -2165 840
rect -2115 920 -2075 930
rect -2115 840 -2105 920
rect -2085 840 -2075 920
rect -2115 830 -2075 840
rect -2025 920 -1985 930
rect -2025 840 -2015 920
rect -1995 840 -1985 920
rect -2025 830 -1985 840
rect -1935 920 -1895 930
rect -1935 840 -1925 920
rect -1905 840 -1895 920
rect -1935 830 -1895 840
rect -1845 920 -1805 930
rect -1845 840 -1835 920
rect -1815 840 -1805 920
rect -1845 830 -1805 840
rect -1755 920 -1715 930
rect -1755 840 -1745 920
rect -1725 840 -1715 920
rect -1755 830 -1715 840
rect -1665 920 -1625 930
rect -1665 840 -1655 920
rect -1635 840 -1625 920
rect -1665 830 -1625 840
rect -1575 920 -1535 930
rect -1575 840 -1565 920
rect -1545 840 -1535 920
rect -1575 830 -1535 840
rect -1485 920 -1445 930
rect -1485 840 -1475 920
rect -1455 840 -1445 920
rect -1485 830 -1445 840
rect -1395 920 -1355 930
rect -1395 840 -1385 920
rect -1365 840 -1355 920
rect -1395 830 -1355 840
rect -1305 920 -1265 930
rect -1305 840 -1295 920
rect -1275 840 -1265 920
rect -1305 830 -1265 840
rect -1215 920 -1175 930
rect -1215 840 -1205 920
rect -1185 840 -1175 920
rect -1215 830 -1175 840
rect -1125 920 -1085 930
rect -1125 840 -1115 920
rect -1095 840 -1085 920
rect -1125 830 -1085 840
rect -1035 920 -995 930
rect -1035 840 -1025 920
rect -1005 840 -995 920
rect -1035 830 -995 840
rect -945 920 -905 930
rect -945 840 -935 920
rect -915 840 -905 920
rect -945 830 -905 840
rect -855 920 -815 930
rect -855 840 -845 920
rect -825 840 -815 920
rect -855 830 -815 840
rect -765 920 -725 930
rect -765 840 -755 920
rect -735 840 -725 920
rect -765 830 -725 840
rect -675 920 -635 930
rect -675 840 -665 920
rect -645 840 -635 920
rect -675 830 -635 840
rect -585 920 -545 930
rect -585 840 -575 920
rect -555 840 -545 920
rect -585 830 -545 840
rect -495 920 -455 930
rect -495 840 -485 920
rect -465 840 -455 920
rect -495 830 -455 840
rect -405 920 -365 930
rect -405 840 -395 920
rect -375 840 -365 920
rect -405 830 -365 840
rect -315 920 -275 930
rect -315 840 -305 920
rect -285 840 -275 920
rect -315 830 -275 840
rect -225 920 -185 930
rect -225 840 -215 920
rect -195 840 -185 920
rect -225 830 -185 840
rect -135 920 -95 930
rect -135 840 -125 920
rect -105 840 -95 920
rect -135 830 -95 840
rect -45 920 -5 930
rect -45 840 -35 920
rect -15 840 -5 920
rect -45 830 -5 840
<< mvndiffc >>
rect -11555 1855 -11535 1935
rect -11465 1855 -11445 1935
rect -11375 1855 -11355 1935
rect -11285 1855 -11265 1935
rect -11195 1855 -11175 1935
rect -11105 1855 -11085 1935
rect -11015 1855 -10995 1935
rect -10925 1855 -10905 1935
rect -10835 1855 -10815 1935
rect -10745 1855 -10725 1935
rect -10655 1855 -10635 1935
rect -10565 1855 -10545 1935
rect -10475 1855 -10455 1935
rect -10385 1855 -10365 1935
rect -10295 1855 -10275 1935
rect -10205 1855 -10185 1935
rect -10115 1855 -10095 1935
rect -10025 1855 -10005 1935
rect -9935 1855 -9915 1935
rect -9845 1855 -9825 1935
rect -9755 1855 -9735 1935
rect -9665 1855 -9645 1935
rect -9575 1855 -9555 1935
rect -9485 1855 -9465 1935
rect -9395 1855 -9375 1935
rect -9305 1855 -9285 1935
rect -9215 1855 -9195 1935
rect -9125 1855 -9105 1935
rect -9035 1855 -9015 1935
rect -8945 1855 -8925 1935
rect -8855 1855 -8835 1935
rect -8765 1855 -8745 1935
rect -8675 1855 -8655 1935
rect -8585 1855 -8565 1935
rect -8495 1855 -8475 1935
rect -8405 1855 -8385 1935
rect -8315 1855 -8295 1935
rect -8225 1855 -8205 1935
rect -8135 1855 -8115 1935
rect -8045 1855 -8025 1935
rect -7955 1855 -7935 1935
rect -7865 1855 -7845 1935
rect -7775 1855 -7755 1935
rect -7685 1855 -7665 1935
rect -7595 1855 -7575 1935
rect -7505 1855 -7485 1935
rect -7415 1855 -7395 1935
rect -7325 1855 -7305 1935
rect -7235 1855 -7215 1935
rect -7145 1855 -7125 1935
rect -7055 1855 -7035 1935
rect -6965 1855 -6945 1935
rect -6875 1855 -6855 1935
rect -6785 1855 -6765 1935
rect -6695 1855 -6675 1935
rect -6605 1855 -6585 1935
rect -6515 1855 -6495 1935
rect -6425 1855 -6405 1935
rect -6335 1855 -6315 1935
rect -6245 1855 -6225 1935
rect -6155 1855 -6135 1935
rect -6065 1855 -6045 1935
rect -5975 1855 -5955 1935
rect -5885 1855 -5865 1935
rect -5795 1855 -5775 1935
rect -5705 1855 -5685 1935
rect -5615 1855 -5595 1935
rect -5525 1855 -5505 1935
rect -5435 1855 -5415 1935
rect -5345 1855 -5325 1935
rect -5255 1855 -5235 1935
rect -5165 1855 -5145 1935
rect -5075 1855 -5055 1935
rect -4985 1855 -4965 1935
rect -4895 1855 -4875 1935
rect -4805 1855 -4785 1935
rect -4715 1855 -4695 1935
rect -4625 1855 -4605 1935
rect -4535 1855 -4515 1935
rect -4445 1855 -4425 1935
rect -4355 1855 -4335 1935
rect -4265 1855 -4245 1935
rect -4175 1855 -4155 1935
rect -4085 1855 -4065 1935
rect -3995 1855 -3975 1935
rect -3905 1855 -3885 1935
rect -3815 1855 -3795 1935
rect -3725 1855 -3705 1935
rect -3635 1855 -3615 1935
rect -3545 1855 -3525 1935
rect -3455 1855 -3435 1935
rect -3365 1855 -3345 1935
rect -3275 1855 -3255 1935
rect -3185 1855 -3165 1935
rect -3095 1855 -3075 1935
rect -3005 1855 -2985 1935
rect -2915 1855 -2895 1935
rect -2825 1855 -2805 1935
rect -2735 1855 -2715 1935
rect -2645 1855 -2625 1935
rect -2555 1855 -2535 1935
rect -2465 1855 -2445 1935
rect -2375 1855 -2355 1935
rect -2285 1855 -2265 1935
rect -2195 1855 -2175 1935
rect -2105 1855 -2085 1935
rect -2015 1855 -1995 1935
rect -1925 1855 -1905 1935
rect -1835 1855 -1815 1935
rect -1745 1855 -1725 1935
rect -1655 1855 -1635 1935
rect -1565 1855 -1545 1935
rect -1475 1855 -1455 1935
rect -1385 1855 -1365 1935
rect -1295 1855 -1275 1935
rect -1205 1855 -1185 1935
rect -1115 1855 -1095 1935
rect -1025 1855 -1005 1935
rect -935 1855 -915 1935
rect -845 1855 -825 1935
rect -755 1855 -735 1935
rect -665 1855 -645 1935
rect -575 1855 -555 1935
rect -485 1855 -465 1935
rect -395 1855 -375 1935
rect -305 1855 -285 1935
rect -215 1855 -195 1935
rect -125 1855 -105 1935
rect -35 1855 -15 1935
rect -11555 60 -11535 140
rect -11465 60 -11445 140
rect -11375 60 -11355 140
rect -11285 60 -11265 140
rect -11195 60 -11175 140
rect -11105 60 -11085 140
rect -11015 60 -10995 140
rect -10925 60 -10905 140
rect -10835 60 -10815 140
rect -10745 60 -10725 140
rect -10655 60 -10635 140
rect -10565 60 -10545 140
rect -10475 60 -10455 140
rect -10385 60 -10365 140
rect -10295 60 -10275 140
rect -10205 60 -10185 140
rect -10115 60 -10095 140
rect -10025 60 -10005 140
rect -9935 60 -9915 140
rect -9845 60 -9825 140
rect -9755 60 -9735 140
rect -9665 60 -9645 140
rect -9575 60 -9555 140
rect -9485 60 -9465 140
rect -9395 60 -9375 140
rect -9305 60 -9285 140
rect -9215 60 -9195 140
rect -9125 60 -9105 140
rect -9035 60 -9015 140
rect -8945 60 -8925 140
rect -8855 60 -8835 140
rect -8765 60 -8745 140
rect -8675 60 -8655 140
rect -8585 60 -8565 140
rect -8495 60 -8475 140
rect -8405 60 -8385 140
rect -8315 60 -8295 140
rect -8225 60 -8205 140
rect -8135 60 -8115 140
rect -8045 60 -8025 140
rect -7955 60 -7935 140
rect -7865 60 -7845 140
rect -7775 60 -7755 140
rect -7685 60 -7665 140
rect -7595 60 -7575 140
rect -7505 60 -7485 140
rect -7415 60 -7395 140
rect -7325 60 -7305 140
rect -7235 60 -7215 140
rect -7145 60 -7125 140
rect -7055 60 -7035 140
rect -6965 60 -6945 140
rect -6875 60 -6855 140
rect -6785 60 -6765 140
rect -6695 60 -6675 140
rect -6605 60 -6585 140
rect -6515 60 -6495 140
rect -6425 60 -6405 140
rect -6335 60 -6315 140
rect -6245 60 -6225 140
rect -6155 60 -6135 140
rect -6065 60 -6045 140
rect -5975 60 -5955 140
rect -5885 60 -5865 140
rect -5795 60 -5775 140
rect -5705 60 -5685 140
rect -5615 60 -5595 140
rect -5525 60 -5505 140
rect -5435 60 -5415 140
rect -5345 60 -5325 140
rect -5255 60 -5235 140
rect -5165 60 -5145 140
rect -5075 60 -5055 140
rect -4985 60 -4965 140
rect -4895 60 -4875 140
rect -4805 60 -4785 140
rect -4715 60 -4695 140
rect -4625 60 -4605 140
rect -4535 60 -4515 140
rect -4445 60 -4425 140
rect -4355 60 -4335 140
rect -4265 60 -4245 140
rect -4175 60 -4155 140
rect -4085 60 -4065 140
rect -3995 60 -3975 140
rect -3905 60 -3885 140
rect -3815 60 -3795 140
rect -3725 60 -3705 140
rect -3635 60 -3615 140
rect -3545 60 -3525 140
rect -3455 60 -3435 140
rect -3365 60 -3345 140
rect -3275 60 -3255 140
rect -3185 60 -3165 140
rect -3095 60 -3075 140
rect -3005 60 -2985 140
rect -2915 60 -2895 140
rect -2825 60 -2805 140
rect -2735 60 -2715 140
rect -2645 60 -2625 140
rect -2555 60 -2535 140
rect -2465 60 -2445 140
rect -2375 60 -2355 140
rect -2285 60 -2265 140
rect -2195 60 -2175 140
rect -2105 60 -2085 140
rect -2015 60 -1995 140
rect -1925 60 -1905 140
rect -1835 60 -1815 140
rect -1745 60 -1725 140
rect -1655 60 -1635 140
rect -1565 60 -1545 140
rect -1475 60 -1455 140
rect -1385 60 -1365 140
rect -1295 60 -1275 140
rect -1205 60 -1185 140
rect -1115 60 -1095 140
rect -1025 60 -1005 140
rect -935 60 -915 140
rect -845 60 -825 140
rect -755 60 -735 140
rect -665 60 -645 140
rect -575 60 -555 140
rect -485 60 -465 140
rect -395 60 -375 140
rect -305 60 -285 140
rect -215 60 -195 140
rect -125 60 -105 140
rect -35 60 -15 140
<< mvpdiffc >>
rect -11555 1075 -11535 1155
rect -11465 1075 -11445 1155
rect -11375 1075 -11355 1155
rect -11285 1075 -11265 1155
rect -11195 1075 -11175 1155
rect -11105 1075 -11085 1155
rect -11015 1075 -10995 1155
rect -10925 1075 -10905 1155
rect -10835 1075 -10815 1155
rect -10745 1075 -10725 1155
rect -10655 1075 -10635 1155
rect -10565 1075 -10545 1155
rect -10475 1075 -10455 1155
rect -10385 1075 -10365 1155
rect -10295 1075 -10275 1155
rect -10205 1075 -10185 1155
rect -10115 1075 -10095 1155
rect -10025 1075 -10005 1155
rect -9935 1075 -9915 1155
rect -9845 1075 -9825 1155
rect -9755 1075 -9735 1155
rect -9665 1075 -9645 1155
rect -9575 1075 -9555 1155
rect -9485 1075 -9465 1155
rect -9395 1075 -9375 1155
rect -9305 1075 -9285 1155
rect -9215 1075 -9195 1155
rect -9125 1075 -9105 1155
rect -9035 1075 -9015 1155
rect -8945 1075 -8925 1155
rect -8855 1075 -8835 1155
rect -8765 1075 -8745 1155
rect -8675 1075 -8655 1155
rect -8585 1075 -8565 1155
rect -8495 1075 -8475 1155
rect -8405 1075 -8385 1155
rect -8315 1075 -8295 1155
rect -8225 1075 -8205 1155
rect -8135 1075 -8115 1155
rect -8045 1075 -8025 1155
rect -7955 1075 -7935 1155
rect -7865 1075 -7845 1155
rect -7775 1075 -7755 1155
rect -7685 1075 -7665 1155
rect -7595 1075 -7575 1155
rect -7505 1075 -7485 1155
rect -7415 1075 -7395 1155
rect -7325 1075 -7305 1155
rect -7235 1075 -7215 1155
rect -7145 1075 -7125 1155
rect -7055 1075 -7035 1155
rect -6965 1075 -6945 1155
rect -6875 1075 -6855 1155
rect -6785 1075 -6765 1155
rect -6695 1075 -6675 1155
rect -6605 1075 -6585 1155
rect -6515 1075 -6495 1155
rect -6425 1075 -6405 1155
rect -6335 1075 -6315 1155
rect -6245 1075 -6225 1155
rect -6155 1075 -6135 1155
rect -6065 1075 -6045 1155
rect -5975 1075 -5955 1155
rect -5885 1075 -5865 1155
rect -5795 1075 -5775 1155
rect -5705 1075 -5685 1155
rect -5615 1075 -5595 1155
rect -5525 1075 -5505 1155
rect -5435 1075 -5415 1155
rect -5345 1075 -5325 1155
rect -5255 1075 -5235 1155
rect -5165 1075 -5145 1155
rect -5075 1075 -5055 1155
rect -4985 1075 -4965 1155
rect -4895 1075 -4875 1155
rect -4805 1075 -4785 1155
rect -4715 1075 -4695 1155
rect -4625 1075 -4605 1155
rect -4535 1075 -4515 1155
rect -4445 1075 -4425 1155
rect -4355 1075 -4335 1155
rect -4265 1075 -4245 1155
rect -4175 1075 -4155 1155
rect -4085 1075 -4065 1155
rect -3995 1075 -3975 1155
rect -3905 1075 -3885 1155
rect -3815 1075 -3795 1155
rect -3725 1075 -3705 1155
rect -3635 1075 -3615 1155
rect -3545 1075 -3525 1155
rect -3455 1075 -3435 1155
rect -3365 1075 -3345 1155
rect -3275 1075 -3255 1155
rect -3185 1075 -3165 1155
rect -3095 1075 -3075 1155
rect -3005 1075 -2985 1155
rect -2915 1075 -2895 1155
rect -2825 1075 -2805 1155
rect -2735 1075 -2715 1155
rect -2645 1075 -2625 1155
rect -2555 1075 -2535 1155
rect -2465 1075 -2445 1155
rect -2375 1075 -2355 1155
rect -2285 1075 -2265 1155
rect -2195 1075 -2175 1155
rect -2105 1075 -2085 1155
rect -2015 1075 -1995 1155
rect -1925 1075 -1905 1155
rect -1835 1075 -1815 1155
rect -1745 1075 -1725 1155
rect -1655 1075 -1635 1155
rect -1565 1075 -1545 1155
rect -1475 1075 -1455 1155
rect -1385 1075 -1365 1155
rect -1295 1075 -1275 1155
rect -1205 1075 -1185 1155
rect -1115 1075 -1095 1155
rect -1025 1075 -1005 1155
rect -935 1075 -915 1155
rect -845 1075 -825 1155
rect -755 1075 -735 1155
rect -665 1075 -645 1155
rect -575 1075 -555 1155
rect -485 1075 -465 1155
rect -395 1075 -375 1155
rect -305 1075 -285 1155
rect -215 1075 -195 1155
rect -125 1075 -105 1155
rect -35 1075 -15 1155
rect -11555 840 -11535 920
rect -11465 840 -11445 920
rect -11375 840 -11355 920
rect -11285 840 -11265 920
rect -11195 840 -11175 920
rect -11105 840 -11085 920
rect -11015 840 -10995 920
rect -10925 840 -10905 920
rect -10835 840 -10815 920
rect -10745 840 -10725 920
rect -10655 840 -10635 920
rect -10565 840 -10545 920
rect -10475 840 -10455 920
rect -10385 840 -10365 920
rect -10295 840 -10275 920
rect -10205 840 -10185 920
rect -10115 840 -10095 920
rect -10025 840 -10005 920
rect -9935 840 -9915 920
rect -9845 840 -9825 920
rect -9755 840 -9735 920
rect -9665 840 -9645 920
rect -9575 840 -9555 920
rect -9485 840 -9465 920
rect -9395 840 -9375 920
rect -9305 840 -9285 920
rect -9215 840 -9195 920
rect -9125 840 -9105 920
rect -9035 840 -9015 920
rect -8945 840 -8925 920
rect -8855 840 -8835 920
rect -8765 840 -8745 920
rect -8675 840 -8655 920
rect -8585 840 -8565 920
rect -8495 840 -8475 920
rect -8405 840 -8385 920
rect -8315 840 -8295 920
rect -8225 840 -8205 920
rect -8135 840 -8115 920
rect -8045 840 -8025 920
rect -7955 840 -7935 920
rect -7865 840 -7845 920
rect -7775 840 -7755 920
rect -7685 840 -7665 920
rect -7595 840 -7575 920
rect -7505 840 -7485 920
rect -7415 840 -7395 920
rect -7325 840 -7305 920
rect -7235 840 -7215 920
rect -7145 840 -7125 920
rect -7055 840 -7035 920
rect -6965 840 -6945 920
rect -6875 840 -6855 920
rect -6785 840 -6765 920
rect -6695 840 -6675 920
rect -6605 840 -6585 920
rect -6515 840 -6495 920
rect -6425 840 -6405 920
rect -6335 840 -6315 920
rect -6245 840 -6225 920
rect -6155 840 -6135 920
rect -6065 840 -6045 920
rect -5975 840 -5955 920
rect -5885 840 -5865 920
rect -5795 840 -5775 920
rect -5705 840 -5685 920
rect -5615 840 -5595 920
rect -5525 840 -5505 920
rect -5435 840 -5415 920
rect -5345 840 -5325 920
rect -5255 840 -5235 920
rect -5165 840 -5145 920
rect -5075 840 -5055 920
rect -4985 840 -4965 920
rect -4895 840 -4875 920
rect -4805 840 -4785 920
rect -4715 840 -4695 920
rect -4625 840 -4605 920
rect -4535 840 -4515 920
rect -4445 840 -4425 920
rect -4355 840 -4335 920
rect -4265 840 -4245 920
rect -4175 840 -4155 920
rect -4085 840 -4065 920
rect -3995 840 -3975 920
rect -3905 840 -3885 920
rect -3815 840 -3795 920
rect -3725 840 -3705 920
rect -3635 840 -3615 920
rect -3545 840 -3525 920
rect -3455 840 -3435 920
rect -3365 840 -3345 920
rect -3275 840 -3255 920
rect -3185 840 -3165 920
rect -3095 840 -3075 920
rect -3005 840 -2985 920
rect -2915 840 -2895 920
rect -2825 840 -2805 920
rect -2735 840 -2715 920
rect -2645 840 -2625 920
rect -2555 840 -2535 920
rect -2465 840 -2445 920
rect -2375 840 -2355 920
rect -2285 840 -2265 920
rect -2195 840 -2175 920
rect -2105 840 -2085 920
rect -2015 840 -1995 920
rect -1925 840 -1905 920
rect -1835 840 -1815 920
rect -1745 840 -1725 920
rect -1655 840 -1635 920
rect -1565 840 -1545 920
rect -1475 840 -1455 920
rect -1385 840 -1365 920
rect -1295 840 -1275 920
rect -1205 840 -1185 920
rect -1115 840 -1095 920
rect -1025 840 -1005 920
rect -935 840 -915 920
rect -845 840 -825 920
rect -755 840 -735 920
rect -665 840 -645 920
rect -575 840 -555 920
rect -485 840 -465 920
rect -395 840 -375 920
rect -305 840 -285 920
rect -215 840 -195 920
rect -125 840 -105 920
rect -35 840 -15 920
<< psubdiff >>
rect -11700 1975 -11510 1995
rect -11490 1975 -11420 1995
rect -11400 1975 -11330 1995
rect -11310 1975 -11240 1995
rect -11220 1975 -11150 1995
rect -11130 1975 -11060 1995
rect -11040 1975 -10970 1995
rect -10950 1975 -10880 1995
rect -10860 1975 -10790 1995
rect -10770 1975 -10700 1995
rect -10680 1975 -10610 1995
rect -10590 1975 -10520 1995
rect -10500 1975 -10430 1995
rect -10410 1975 -10340 1995
rect -10320 1975 -10250 1995
rect -10230 1975 -10160 1995
rect -10140 1975 -10070 1995
rect -10050 1975 -9980 1995
rect -9960 1975 -9890 1995
rect -9870 1975 -9800 1995
rect -9780 1975 -9710 1995
rect -9690 1975 -9620 1995
rect -9600 1975 -9530 1995
rect -9510 1975 -9440 1995
rect -9420 1975 -9350 1995
rect -9330 1975 -9260 1995
rect -9240 1975 -9170 1995
rect -9150 1975 -9080 1995
rect -9060 1975 -8990 1995
rect -8970 1975 -8900 1995
rect -8880 1975 -8810 1995
rect -8790 1975 -8720 1995
rect -8700 1975 -8630 1995
rect -8610 1975 -8540 1995
rect -8520 1975 -8450 1995
rect -8430 1975 -8360 1995
rect -8340 1975 -8270 1995
rect -8250 1975 -8180 1995
rect -8160 1975 -8090 1995
rect -8070 1975 -8000 1995
rect -7980 1975 -7910 1995
rect -7890 1975 -7820 1995
rect -7800 1975 -7730 1995
rect -7710 1975 -7640 1995
rect -7620 1975 -7550 1995
rect -7530 1975 -7460 1995
rect -7440 1975 -7370 1995
rect -7350 1975 -7280 1995
rect -7260 1975 -7190 1995
rect -7170 1975 -7100 1995
rect -7080 1975 -7010 1995
rect -6990 1975 -6920 1995
rect -6900 1975 -6830 1995
rect -6810 1975 -6740 1995
rect -6720 1975 -6650 1995
rect -6630 1975 -6560 1995
rect -6540 1975 -6470 1995
rect -6450 1975 -6380 1995
rect -6360 1975 -6290 1995
rect -6270 1975 -6200 1995
rect -6180 1975 -6110 1995
rect -6090 1975 -6020 1995
rect -6000 1975 -5930 1995
rect -5910 1975 -5840 1995
rect -5820 1975 -5750 1995
rect -5730 1975 -5660 1995
rect -5640 1975 -5570 1995
rect -5550 1975 -5480 1995
rect -5460 1975 -5390 1995
rect -5370 1975 -5300 1995
rect -5280 1975 -5210 1995
rect -5190 1975 -5120 1995
rect -5100 1975 -5030 1995
rect -5010 1975 -4940 1995
rect -4920 1975 -4850 1995
rect -4830 1975 -4760 1995
rect -4740 1975 -4670 1995
rect -4650 1975 -4580 1995
rect -4560 1975 -4490 1995
rect -4470 1975 -4400 1995
rect -4380 1975 -4310 1995
rect -4290 1975 -4220 1995
rect -4200 1975 -4130 1995
rect -4110 1975 -4040 1995
rect -4020 1975 -3950 1995
rect -3930 1975 -3860 1995
rect -3840 1975 -3770 1995
rect -3750 1975 -3680 1995
rect -3660 1975 -3590 1995
rect -3570 1975 -3500 1995
rect -3480 1975 -3410 1995
rect -3390 1975 -3320 1995
rect -3300 1975 -3230 1995
rect -3210 1975 -3140 1995
rect -3120 1975 -3050 1995
rect -3030 1975 -2960 1995
rect -2940 1975 -2870 1995
rect -2850 1975 -2780 1995
rect -2760 1975 -2690 1995
rect -2670 1975 -2600 1995
rect -2580 1975 -2510 1995
rect -2490 1975 -2420 1995
rect -2400 1975 -2330 1995
rect -2310 1975 -2240 1995
rect -2220 1975 -2150 1995
rect -2130 1975 -2060 1995
rect -2040 1975 -1970 1995
rect -1950 1975 -1880 1995
rect -1860 1975 -1790 1995
rect -1770 1975 -1700 1995
rect -1680 1975 -1610 1995
rect -1590 1975 -1520 1995
rect -1500 1975 -1430 1995
rect -1410 1975 -1340 1995
rect -1320 1975 -1250 1995
rect -1230 1975 -1160 1995
rect -1140 1975 -1070 1995
rect -1050 1975 -980 1995
rect -960 1975 -890 1995
rect -870 1975 -800 1995
rect -780 1975 -710 1995
rect -690 1975 -620 1995
rect -600 1975 -530 1995
rect -510 1975 -440 1995
rect -420 1975 -350 1995
rect -330 1975 -260 1995
rect -240 1975 -170 1995
rect -150 1975 -80 1995
rect -60 1975 130 1995
rect -11690 1775 -11670 1975
rect 100 1775 120 1975
rect -11690 1755 -11510 1775
rect -11490 1755 -11420 1775
rect -11400 1755 -11330 1775
rect -11310 1755 -11240 1775
rect -11220 1755 -11150 1775
rect -11130 1755 -11060 1775
rect -11040 1755 -10970 1775
rect -10950 1755 -10880 1775
rect -10860 1755 -10790 1775
rect -10770 1755 -10700 1775
rect -10680 1755 -10610 1775
rect -10590 1755 -10520 1775
rect -10500 1755 -10430 1775
rect -10410 1755 -10340 1775
rect -10320 1755 -10250 1775
rect -10230 1755 -10160 1775
rect -10140 1755 -10070 1775
rect -10050 1755 -9980 1775
rect -9960 1755 -9890 1775
rect -9870 1755 -9800 1775
rect -9780 1755 -9710 1775
rect -9690 1755 -9620 1775
rect -9600 1755 -9530 1775
rect -9510 1755 -9440 1775
rect -9420 1755 -9350 1775
rect -9330 1755 -9260 1775
rect -9240 1755 -9170 1775
rect -9150 1755 -9080 1775
rect -9060 1755 -8990 1775
rect -8970 1755 -8900 1775
rect -8880 1755 -8810 1775
rect -8790 1755 -8720 1775
rect -8700 1755 -8630 1775
rect -8610 1755 -8540 1775
rect -8520 1755 -8450 1775
rect -8430 1755 -8360 1775
rect -8340 1755 -8270 1775
rect -8250 1755 -8180 1775
rect -8160 1755 -8090 1775
rect -8070 1755 -8000 1775
rect -7980 1755 -7910 1775
rect -7890 1755 -7820 1775
rect -7800 1755 -7730 1775
rect -7710 1755 -7640 1775
rect -7620 1755 -7550 1775
rect -7530 1755 -7460 1775
rect -7440 1755 -7370 1775
rect -7350 1755 -7280 1775
rect -7260 1755 -7190 1775
rect -7170 1755 -7100 1775
rect -7080 1755 -7010 1775
rect -6990 1755 -6920 1775
rect -6900 1755 -6830 1775
rect -6810 1755 -6740 1775
rect -6720 1755 -6650 1775
rect -6630 1755 -6560 1775
rect -6540 1755 -6470 1775
rect -6450 1755 -6380 1775
rect -6360 1755 -6290 1775
rect -6270 1755 -6200 1775
rect -6180 1755 -6110 1775
rect -6090 1755 -6020 1775
rect -6000 1755 -5930 1775
rect -5910 1755 -5840 1775
rect -5820 1755 -5750 1775
rect -5730 1755 -5660 1775
rect -5640 1755 -5570 1775
rect -5550 1755 -5480 1775
rect -5460 1755 -5390 1775
rect -5370 1755 -5300 1775
rect -5280 1755 -5210 1775
rect -5190 1755 -5120 1775
rect -5100 1755 -5030 1775
rect -5010 1755 -4940 1775
rect -4920 1755 -4850 1775
rect -4830 1755 -4760 1775
rect -4740 1755 -4670 1775
rect -4650 1755 -4580 1775
rect -4560 1755 -4490 1775
rect -4470 1755 -4400 1775
rect -4380 1755 -4310 1775
rect -4290 1755 -4220 1775
rect -4200 1755 -4130 1775
rect -4110 1755 -4040 1775
rect -4020 1755 -3950 1775
rect -3930 1755 -3860 1775
rect -3840 1755 -3770 1775
rect -3750 1755 -3680 1775
rect -3660 1755 -3590 1775
rect -3570 1755 -3500 1775
rect -3480 1755 -3410 1775
rect -3390 1755 -3320 1775
rect -3300 1755 -3230 1775
rect -3210 1755 -3140 1775
rect -3120 1755 -3050 1775
rect -3030 1755 -2960 1775
rect -2940 1755 -2870 1775
rect -2850 1755 -2780 1775
rect -2760 1755 -2690 1775
rect -2670 1755 -2600 1775
rect -2580 1755 -2510 1775
rect -2490 1755 -2420 1775
rect -2400 1755 -2330 1775
rect -2310 1755 -2240 1775
rect -2220 1755 -2150 1775
rect -2130 1755 -2060 1775
rect -2040 1755 -1970 1775
rect -1950 1755 -1880 1775
rect -1860 1755 -1790 1775
rect -1770 1755 -1700 1775
rect -1680 1755 -1610 1775
rect -1590 1755 -1520 1775
rect -1500 1755 -1430 1775
rect -1410 1755 -1340 1775
rect -1320 1755 -1250 1775
rect -1230 1755 -1160 1775
rect -1140 1755 -1070 1775
rect -1050 1755 -980 1775
rect -960 1755 -890 1775
rect -870 1755 -800 1775
rect -780 1755 -710 1775
rect -690 1755 -620 1775
rect -600 1755 -530 1775
rect -510 1755 -440 1775
rect -420 1755 -350 1775
rect -330 1755 -260 1775
rect -240 1755 -170 1775
rect -150 1755 -80 1775
rect -60 1755 120 1775
rect -11690 1315 -11510 1335
rect -11490 1315 -11420 1335
rect -11400 1315 -11330 1335
rect -11310 1315 -11240 1335
rect -11220 1315 -11150 1335
rect -11130 1315 -11060 1335
rect -11040 1315 -10970 1335
rect -10950 1315 -10880 1335
rect -10860 1315 -10790 1335
rect -10770 1315 -10700 1335
rect -10680 1315 -10610 1335
rect -10590 1315 -10520 1335
rect -10500 1315 -10430 1335
rect -10410 1315 -10340 1335
rect -10320 1315 -10250 1335
rect -10230 1315 -10160 1335
rect -10140 1315 -10070 1335
rect -10050 1315 -9980 1335
rect -9960 1315 -9890 1335
rect -9870 1315 -9800 1335
rect -9780 1315 -9710 1335
rect -9690 1315 -9620 1335
rect -9600 1315 -9530 1335
rect -9510 1315 -9440 1335
rect -9420 1315 -9350 1335
rect -9330 1315 -9260 1335
rect -9240 1315 -9170 1335
rect -9150 1315 -9080 1335
rect -9060 1315 -8990 1335
rect -8970 1315 -8900 1335
rect -8880 1315 -8810 1335
rect -8790 1315 -8720 1335
rect -8700 1315 -8630 1335
rect -8610 1315 -8540 1335
rect -8520 1315 -8450 1335
rect -8430 1315 -8360 1335
rect -8340 1315 -8270 1335
rect -8250 1315 -8180 1335
rect -8160 1315 -8090 1335
rect -8070 1315 -8000 1335
rect -7980 1315 -7910 1335
rect -7890 1315 -7820 1335
rect -7800 1315 -7730 1335
rect -7710 1315 -7640 1335
rect -7620 1315 -7550 1335
rect -7530 1315 -7460 1335
rect -7440 1315 -7370 1335
rect -7350 1315 -7280 1335
rect -7260 1315 -7190 1335
rect -7170 1315 -7100 1335
rect -7080 1315 -7010 1335
rect -6990 1315 -6920 1335
rect -6900 1315 -6830 1335
rect -6810 1315 -6740 1335
rect -6720 1315 -6650 1335
rect -6630 1315 -6560 1335
rect -6540 1315 -6470 1335
rect -6450 1315 -6380 1335
rect -6360 1315 -6290 1335
rect -6270 1315 -6200 1335
rect -6180 1315 -6110 1335
rect -6090 1315 -6020 1335
rect -6000 1315 -5930 1335
rect -5910 1315 -5840 1335
rect -5820 1315 -5750 1335
rect -5730 1315 -5660 1335
rect -5640 1315 -5570 1335
rect -5550 1315 -5480 1335
rect -5460 1315 -5390 1335
rect -5370 1315 -5300 1335
rect -5280 1315 -5210 1335
rect -5190 1315 -5120 1335
rect -5100 1315 -5030 1335
rect -5010 1315 -4940 1335
rect -4920 1315 -4850 1335
rect -4830 1315 -4760 1335
rect -4740 1315 -4670 1335
rect -4650 1315 -4580 1335
rect -4560 1315 -4490 1335
rect -4470 1315 -4400 1335
rect -4380 1315 -4310 1335
rect -4290 1315 -4220 1335
rect -4200 1315 -4130 1335
rect -4110 1315 -4040 1335
rect -4020 1315 -3950 1335
rect -3930 1315 -3860 1335
rect -3840 1315 -3770 1335
rect -3750 1315 -3680 1335
rect -3660 1315 -3590 1335
rect -3570 1315 -3500 1335
rect -3480 1315 -3410 1335
rect -3390 1315 -3320 1335
rect -3300 1315 -3230 1335
rect -3210 1315 -3140 1335
rect -3120 1315 -3050 1335
rect -3030 1315 -2960 1335
rect -2940 1315 -2870 1335
rect -2850 1315 -2780 1335
rect -2760 1315 -2690 1335
rect -2670 1315 -2600 1335
rect -2580 1315 -2510 1335
rect -2490 1315 -2420 1335
rect -2400 1315 -2330 1335
rect -2310 1315 -2240 1335
rect -2220 1315 -2150 1335
rect -2130 1315 -2060 1335
rect -2040 1315 -1970 1335
rect -1950 1315 -1880 1335
rect -1860 1315 -1790 1335
rect -1770 1315 -1700 1335
rect -1680 1315 -1610 1335
rect -1590 1315 -1520 1335
rect -1500 1315 -1430 1335
rect -1410 1315 -1340 1335
rect -1320 1315 -1250 1335
rect -1230 1315 -1160 1335
rect -1140 1315 -1070 1335
rect -1050 1315 -980 1335
rect -960 1315 -890 1335
rect -870 1315 -800 1335
rect -780 1315 -710 1335
rect -690 1315 -620 1335
rect -600 1315 -530 1335
rect -510 1315 -440 1335
rect -420 1315 -350 1335
rect -330 1315 -260 1335
rect -240 1315 -170 1335
rect -150 1315 -80 1335
rect -60 1315 120 1335
rect -11690 680 -11670 1315
rect 100 680 120 1315
rect -11690 660 -11510 680
rect -11490 660 -11420 680
rect -11400 660 -11330 680
rect -11310 660 -11240 680
rect -11220 660 -11150 680
rect -11130 660 -11060 680
rect -11040 660 -10970 680
rect -10950 660 -10880 680
rect -10860 660 -10790 680
rect -10770 660 -10700 680
rect -10680 660 -10610 680
rect -10590 660 -10520 680
rect -10500 660 -10430 680
rect -10410 660 -10340 680
rect -10320 660 -10250 680
rect -10230 660 -10160 680
rect -10140 660 -10070 680
rect -10050 660 -9980 680
rect -9960 660 -9890 680
rect -9870 660 -9800 680
rect -9780 660 -9710 680
rect -9690 660 -9620 680
rect -9600 660 -9530 680
rect -9510 660 -9440 680
rect -9420 660 -9350 680
rect -9330 660 -9260 680
rect -9240 660 -9170 680
rect -9150 660 -9080 680
rect -9060 660 -8990 680
rect -8970 660 -8900 680
rect -8880 660 -8810 680
rect -8790 660 -8720 680
rect -8700 660 -8630 680
rect -8610 660 -8540 680
rect -8520 660 -8450 680
rect -8430 660 -8360 680
rect -8340 660 -8270 680
rect -8250 660 -8180 680
rect -8160 660 -8090 680
rect -8070 660 -8000 680
rect -7980 660 -7910 680
rect -7890 660 -7820 680
rect -7800 660 -7730 680
rect -7710 660 -7640 680
rect -7620 660 -7550 680
rect -7530 660 -7460 680
rect -7440 660 -7370 680
rect -7350 660 -7280 680
rect -7260 660 -7190 680
rect -7170 660 -7100 680
rect -7080 660 -7010 680
rect -6990 660 -6920 680
rect -6900 660 -6830 680
rect -6810 660 -6740 680
rect -6720 660 -6650 680
rect -6630 660 -6560 680
rect -6540 660 -6470 680
rect -6450 660 -6380 680
rect -6360 660 -6290 680
rect -6270 660 -6200 680
rect -6180 660 -6110 680
rect -6090 660 -6020 680
rect -6000 660 -5930 680
rect -5910 660 -5840 680
rect -5820 660 -5750 680
rect -5730 660 -5660 680
rect -5640 660 -5570 680
rect -5550 660 -5480 680
rect -5460 660 -5390 680
rect -5370 660 -5300 680
rect -5280 660 -5210 680
rect -5190 660 -5120 680
rect -5100 660 -5030 680
rect -5010 660 -4940 680
rect -4920 660 -4850 680
rect -4830 660 -4760 680
rect -4740 660 -4670 680
rect -4650 660 -4580 680
rect -4560 660 -4490 680
rect -4470 660 -4400 680
rect -4380 660 -4310 680
rect -4290 660 -4220 680
rect -4200 660 -4130 680
rect -4110 660 -4040 680
rect -4020 660 -3950 680
rect -3930 660 -3860 680
rect -3840 660 -3770 680
rect -3750 660 -3680 680
rect -3660 660 -3590 680
rect -3570 660 -3500 680
rect -3480 660 -3410 680
rect -3390 660 -3320 680
rect -3300 660 -3230 680
rect -3210 660 -3140 680
rect -3120 660 -3050 680
rect -3030 660 -2960 680
rect -2940 660 -2870 680
rect -2850 660 -2780 680
rect -2760 660 -2690 680
rect -2670 660 -2600 680
rect -2580 660 -2510 680
rect -2490 660 -2420 680
rect -2400 660 -2330 680
rect -2310 660 -2240 680
rect -2220 660 -2150 680
rect -2130 660 -2060 680
rect -2040 660 -1970 680
rect -1950 660 -1880 680
rect -1860 660 -1790 680
rect -1770 660 -1700 680
rect -1680 660 -1610 680
rect -1590 660 -1520 680
rect -1500 660 -1430 680
rect -1410 660 -1340 680
rect -1320 660 -1250 680
rect -1230 660 -1160 680
rect -1140 660 -1070 680
rect -1050 660 -980 680
rect -960 660 -890 680
rect -870 660 -800 680
rect -780 660 -710 680
rect -690 660 -620 680
rect -600 660 -530 680
rect -510 660 -440 680
rect -420 660 -350 680
rect -330 660 -260 680
rect -240 660 -170 680
rect -150 660 -80 680
rect -60 660 120 680
rect -11690 220 -11510 240
rect -11490 220 -11420 240
rect -11400 220 -11330 240
rect -11310 220 -11240 240
rect -11220 220 -11150 240
rect -11130 220 -11060 240
rect -11040 220 -10970 240
rect -10950 220 -10880 240
rect -10860 220 -10790 240
rect -10770 220 -10700 240
rect -10680 220 -10610 240
rect -10590 220 -10520 240
rect -10500 220 -10430 240
rect -10410 220 -10340 240
rect -10320 220 -10250 240
rect -10230 220 -10160 240
rect -10140 220 -10070 240
rect -10050 220 -9980 240
rect -9960 220 -9890 240
rect -9870 220 -9800 240
rect -9780 220 -9710 240
rect -9690 220 -9620 240
rect -9600 220 -9530 240
rect -9510 220 -9440 240
rect -9420 220 -9350 240
rect -9330 220 -9260 240
rect -9240 220 -9170 240
rect -9150 220 -9080 240
rect -9060 220 -8990 240
rect -8970 220 -8900 240
rect -8880 220 -8810 240
rect -8790 220 -8720 240
rect -8700 220 -8630 240
rect -8610 220 -8540 240
rect -8520 220 -8450 240
rect -8430 220 -8360 240
rect -8340 220 -8270 240
rect -8250 220 -8180 240
rect -8160 220 -8090 240
rect -8070 220 -8000 240
rect -7980 220 -7910 240
rect -7890 220 -7820 240
rect -7800 220 -7730 240
rect -7710 220 -7640 240
rect -7620 220 -7550 240
rect -7530 220 -7460 240
rect -7440 220 -7370 240
rect -7350 220 -7280 240
rect -7260 220 -7190 240
rect -7170 220 -7100 240
rect -7080 220 -7010 240
rect -6990 220 -6920 240
rect -6900 220 -6830 240
rect -6810 220 -6740 240
rect -6720 220 -6650 240
rect -6630 220 -6560 240
rect -6540 220 -6470 240
rect -6450 220 -6380 240
rect -6360 220 -6290 240
rect -6270 220 -6200 240
rect -6180 220 -6110 240
rect -6090 220 -6020 240
rect -6000 220 -5930 240
rect -5910 220 -5840 240
rect -5820 220 -5750 240
rect -5730 220 -5660 240
rect -5640 220 -5570 240
rect -5550 220 -5480 240
rect -5460 220 -5390 240
rect -5370 220 -5300 240
rect -5280 220 -5210 240
rect -5190 220 -5120 240
rect -5100 220 -5030 240
rect -5010 220 -4940 240
rect -4920 220 -4850 240
rect -4830 220 -4760 240
rect -4740 220 -4670 240
rect -4650 220 -4580 240
rect -4560 220 -4490 240
rect -4470 220 -4400 240
rect -4380 220 -4310 240
rect -4290 220 -4220 240
rect -4200 220 -4130 240
rect -4110 220 -4040 240
rect -4020 220 -3950 240
rect -3930 220 -3860 240
rect -3840 220 -3770 240
rect -3750 220 -3680 240
rect -3660 220 -3590 240
rect -3570 220 -3500 240
rect -3480 220 -3410 240
rect -3390 220 -3320 240
rect -3300 220 -3230 240
rect -3210 220 -3140 240
rect -3120 220 -3050 240
rect -3030 220 -2960 240
rect -2940 220 -2870 240
rect -2850 220 -2780 240
rect -2760 220 -2690 240
rect -2670 220 -2600 240
rect -2580 220 -2510 240
rect -2490 220 -2420 240
rect -2400 220 -2330 240
rect -2310 220 -2240 240
rect -2220 220 -2150 240
rect -2130 220 -2060 240
rect -2040 220 -1970 240
rect -1950 220 -1880 240
rect -1860 220 -1790 240
rect -1770 220 -1700 240
rect -1680 220 -1610 240
rect -1590 220 -1520 240
rect -1500 220 -1430 240
rect -1410 220 -1340 240
rect -1320 220 -1250 240
rect -1230 220 -1160 240
rect -1140 220 -1070 240
rect -1050 220 -980 240
rect -960 220 -890 240
rect -870 220 -800 240
rect -780 220 -710 240
rect -690 220 -620 240
rect -600 220 -530 240
rect -510 220 -440 240
rect -420 220 -350 240
rect -330 220 -260 240
rect -240 220 -170 240
rect -150 220 -80 240
rect -60 220 120 240
rect -11690 20 -11670 220
rect 100 20 120 220
rect -11700 0 -11510 20
rect -11490 0 -11420 20
rect -11400 0 -11330 20
rect -11310 0 -11240 20
rect -11220 0 -11150 20
rect -11130 0 -11060 20
rect -11040 0 -10970 20
rect -10950 0 -10880 20
rect -10860 0 -10790 20
rect -10770 0 -10700 20
rect -10680 0 -10610 20
rect -10590 0 -10520 20
rect -10500 0 -10430 20
rect -10410 0 -10340 20
rect -10320 0 -10250 20
rect -10230 0 -10160 20
rect -10140 0 -10070 20
rect -10050 0 -9980 20
rect -9960 0 -9890 20
rect -9870 0 -9800 20
rect -9780 0 -9710 20
rect -9690 0 -9620 20
rect -9600 0 -9530 20
rect -9510 0 -9440 20
rect -9420 0 -9350 20
rect -9330 0 -9260 20
rect -9240 0 -9170 20
rect -9150 0 -9080 20
rect -9060 0 -8990 20
rect -8970 0 -8900 20
rect -8880 0 -8810 20
rect -8790 0 -8720 20
rect -8700 0 -8630 20
rect -8610 0 -8540 20
rect -8520 0 -8450 20
rect -8430 0 -8360 20
rect -8340 0 -8270 20
rect -8250 0 -8180 20
rect -8160 0 -8090 20
rect -8070 0 -8000 20
rect -7980 0 -7910 20
rect -7890 0 -7820 20
rect -7800 0 -7730 20
rect -7710 0 -7640 20
rect -7620 0 -7550 20
rect -7530 0 -7460 20
rect -7440 0 -7370 20
rect -7350 0 -7280 20
rect -7260 0 -7190 20
rect -7170 0 -7100 20
rect -7080 0 -7010 20
rect -6990 0 -6920 20
rect -6900 0 -6830 20
rect -6810 0 -6740 20
rect -6720 0 -6650 20
rect -6630 0 -6560 20
rect -6540 0 -6470 20
rect -6450 0 -6380 20
rect -6360 0 -6290 20
rect -6270 0 -6200 20
rect -6180 0 -6110 20
rect -6090 0 -6020 20
rect -6000 0 -5930 20
rect -5910 0 -5840 20
rect -5820 0 -5750 20
rect -5730 0 -5660 20
rect -5640 0 -5570 20
rect -5550 0 -5480 20
rect -5460 0 -5390 20
rect -5370 0 -5300 20
rect -5280 0 -5210 20
rect -5190 0 -5120 20
rect -5100 0 -5030 20
rect -5010 0 -4940 20
rect -4920 0 -4850 20
rect -4830 0 -4760 20
rect -4740 0 -4670 20
rect -4650 0 -4580 20
rect -4560 0 -4490 20
rect -4470 0 -4400 20
rect -4380 0 -4310 20
rect -4290 0 -4220 20
rect -4200 0 -4130 20
rect -4110 0 -4040 20
rect -4020 0 -3950 20
rect -3930 0 -3860 20
rect -3840 0 -3770 20
rect -3750 0 -3680 20
rect -3660 0 -3590 20
rect -3570 0 -3500 20
rect -3480 0 -3410 20
rect -3390 0 -3320 20
rect -3300 0 -3230 20
rect -3210 0 -3140 20
rect -3120 0 -3050 20
rect -3030 0 -2960 20
rect -2940 0 -2870 20
rect -2850 0 -2780 20
rect -2760 0 -2690 20
rect -2670 0 -2600 20
rect -2580 0 -2510 20
rect -2490 0 -2420 20
rect -2400 0 -2330 20
rect -2310 0 -2240 20
rect -2220 0 -2150 20
rect -2130 0 -2060 20
rect -2040 0 -1970 20
rect -1950 0 -1880 20
rect -1860 0 -1790 20
rect -1770 0 -1700 20
rect -1680 0 -1610 20
rect -1590 0 -1520 20
rect -1500 0 -1430 20
rect -1410 0 -1340 20
rect -1320 0 -1250 20
rect -1230 0 -1160 20
rect -1140 0 -1070 20
rect -1050 0 -980 20
rect -960 0 -890 20
rect -870 0 -800 20
rect -780 0 -710 20
rect -690 0 -620 20
rect -600 0 -530 20
rect -510 0 -440 20
rect -420 0 -350 20
rect -330 0 -260 20
rect -240 0 -170 20
rect -150 0 -80 20
rect -60 0 130 20
<< nsubdiff >>
rect -11615 1235 -11510 1255
rect -11490 1235 -11420 1255
rect -11400 1235 -11330 1255
rect -11310 1235 -11240 1255
rect -11220 1235 -11150 1255
rect -11130 1235 -11060 1255
rect -11040 1235 -10970 1255
rect -10950 1235 -10880 1255
rect -10860 1235 -10790 1255
rect -10770 1235 -10700 1255
rect -10680 1235 -10610 1255
rect -10590 1235 -10520 1255
rect -10500 1235 -10430 1255
rect -10410 1235 -10340 1255
rect -10320 1235 -10250 1255
rect -10230 1235 -10160 1255
rect -10140 1235 -10070 1255
rect -10050 1235 -9980 1255
rect -9960 1235 -9890 1255
rect -9870 1235 -9800 1255
rect -9780 1235 -9710 1255
rect -9690 1235 -9620 1255
rect -9600 1235 -9530 1255
rect -9510 1235 -9440 1255
rect -9420 1235 -9350 1255
rect -9330 1235 -9260 1255
rect -9240 1235 -9170 1255
rect -9150 1235 -9080 1255
rect -9060 1235 -8990 1255
rect -8970 1235 -8900 1255
rect -8880 1235 -8810 1255
rect -8790 1235 -8720 1255
rect -8700 1235 -8630 1255
rect -8610 1235 -8540 1255
rect -8520 1235 -8450 1255
rect -8430 1235 -8360 1255
rect -8340 1235 -8270 1255
rect -8250 1235 -8180 1255
rect -8160 1235 -8090 1255
rect -8070 1235 -8000 1255
rect -7980 1235 -7910 1255
rect -7890 1235 -7820 1255
rect -7800 1235 -7730 1255
rect -7710 1235 -7640 1255
rect -7620 1235 -7550 1255
rect -7530 1235 -7460 1255
rect -7440 1235 -7370 1255
rect -7350 1235 -7280 1255
rect -7260 1235 -7190 1255
rect -7170 1235 -7100 1255
rect -7080 1235 -7010 1255
rect -6990 1235 -6920 1255
rect -6900 1235 -6830 1255
rect -6810 1235 -6740 1255
rect -6720 1235 -6650 1255
rect -6630 1235 -6560 1255
rect -6540 1235 -6470 1255
rect -6450 1235 -6380 1255
rect -6360 1235 -6290 1255
rect -6270 1235 -6200 1255
rect -6180 1235 -6110 1255
rect -6090 1235 -6020 1255
rect -6000 1235 -5930 1255
rect -5910 1235 -5840 1255
rect -5820 1235 -5750 1255
rect -5730 1235 -5660 1255
rect -5640 1235 -5570 1255
rect -5550 1235 -5480 1255
rect -5460 1235 -5390 1255
rect -5370 1235 -5300 1255
rect -5280 1235 -5210 1255
rect -5190 1235 -5120 1255
rect -5100 1235 -5030 1255
rect -5010 1235 -4940 1255
rect -4920 1235 -4850 1255
rect -4830 1235 -4760 1255
rect -4740 1235 -4670 1255
rect -4650 1235 -4580 1255
rect -4560 1235 -4490 1255
rect -4470 1235 -4400 1255
rect -4380 1235 -4310 1255
rect -4290 1235 -4220 1255
rect -4200 1235 -4130 1255
rect -4110 1235 -4040 1255
rect -4020 1235 -3950 1255
rect -3930 1235 -3860 1255
rect -3840 1235 -3770 1255
rect -3750 1235 -3680 1255
rect -3660 1235 -3590 1255
rect -3570 1235 -3500 1255
rect -3480 1235 -3410 1255
rect -3390 1235 -3320 1255
rect -3300 1235 -3230 1255
rect -3210 1235 -3140 1255
rect -3120 1235 -3050 1255
rect -3030 1235 -2960 1255
rect -2940 1235 -2870 1255
rect -2850 1235 -2780 1255
rect -2760 1235 -2690 1255
rect -2670 1235 -2600 1255
rect -2580 1235 -2510 1255
rect -2490 1235 -2420 1255
rect -2400 1235 -2330 1255
rect -2310 1235 -2240 1255
rect -2220 1235 -2150 1255
rect -2130 1235 -2060 1255
rect -2040 1235 -1970 1255
rect -1950 1235 -1880 1255
rect -1860 1235 -1790 1255
rect -1770 1235 -1700 1255
rect -1680 1235 -1610 1255
rect -1590 1235 -1520 1255
rect -1500 1235 -1430 1255
rect -1410 1235 -1340 1255
rect -1320 1235 -1250 1255
rect -1230 1235 -1160 1255
rect -1140 1235 -1070 1255
rect -1050 1235 -980 1255
rect -960 1235 -890 1255
rect -870 1235 -800 1255
rect -780 1235 -710 1255
rect -690 1235 -620 1255
rect -600 1235 -530 1255
rect -510 1235 -440 1255
rect -420 1235 -350 1255
rect -330 1235 -260 1255
rect -240 1235 -170 1255
rect -150 1235 -80 1255
rect -60 1235 45 1255
rect -11615 1035 -11595 1235
rect 25 1035 45 1235
rect -11615 1015 -11510 1035
rect -11490 1015 -11420 1035
rect -11400 1015 -11330 1035
rect -11310 1015 -11240 1035
rect -11220 1015 -11150 1035
rect -11130 1015 -11060 1035
rect -11040 1015 -10970 1035
rect -10950 1015 -10880 1035
rect -10860 1015 -10790 1035
rect -10770 1015 -10700 1035
rect -10680 1015 -10610 1035
rect -10590 1015 -10520 1035
rect -10500 1015 -10430 1035
rect -10410 1015 -10340 1035
rect -10320 1015 -10250 1035
rect -10230 1015 -10160 1035
rect -10140 1015 -10070 1035
rect -10050 1015 -9980 1035
rect -9960 1015 -9890 1035
rect -9870 1015 -9800 1035
rect -9780 1015 -9710 1035
rect -9690 1015 -9620 1035
rect -9600 1015 -9530 1035
rect -9510 1015 -9440 1035
rect -9420 1015 -9350 1035
rect -9330 1015 -9260 1035
rect -9240 1015 -9170 1035
rect -9150 1015 -9080 1035
rect -9060 1015 -8990 1035
rect -8970 1015 -8900 1035
rect -8880 1015 -8810 1035
rect -8790 1015 -8720 1035
rect -8700 1015 -8630 1035
rect -8610 1015 -8540 1035
rect -8520 1015 -8450 1035
rect -8430 1015 -8360 1035
rect -8340 1015 -8270 1035
rect -8250 1015 -8180 1035
rect -8160 1015 -8090 1035
rect -8070 1015 -8000 1035
rect -7980 1015 -7910 1035
rect -7890 1015 -7820 1035
rect -7800 1015 -7730 1035
rect -7710 1015 -7640 1035
rect -7620 1015 -7550 1035
rect -7530 1015 -7460 1035
rect -7440 1015 -7370 1035
rect -7350 1015 -7280 1035
rect -7260 1015 -7190 1035
rect -7170 1015 -7100 1035
rect -7080 1015 -7010 1035
rect -6990 1015 -6920 1035
rect -6900 1015 -6830 1035
rect -6810 1015 -6740 1035
rect -6720 1015 -6650 1035
rect -6630 1015 -6560 1035
rect -6540 1015 -6470 1035
rect -6450 1015 -6380 1035
rect -6360 1015 -6290 1035
rect -6270 1015 -6200 1035
rect -6180 1015 -6110 1035
rect -6090 1015 -6020 1035
rect -6000 1015 -5930 1035
rect -5910 1015 -5840 1035
rect -5820 1015 -5750 1035
rect -5730 1015 -5660 1035
rect -5640 1015 -5570 1035
rect -5550 1015 -5480 1035
rect -5460 1015 -5390 1035
rect -5370 1015 -5300 1035
rect -5280 1015 -5210 1035
rect -5190 1015 -5120 1035
rect -5100 1015 -5030 1035
rect -5010 1015 -4940 1035
rect -4920 1015 -4850 1035
rect -4830 1015 -4760 1035
rect -4740 1015 -4670 1035
rect -4650 1015 -4580 1035
rect -4560 1015 -4490 1035
rect -4470 1015 -4400 1035
rect -4380 1015 -4310 1035
rect -4290 1015 -4220 1035
rect -4200 1015 -4130 1035
rect -4110 1015 -4040 1035
rect -4020 1015 -3950 1035
rect -3930 1015 -3860 1035
rect -3840 1015 -3770 1035
rect -3750 1015 -3680 1035
rect -3660 1015 -3590 1035
rect -3570 1015 -3500 1035
rect -3480 1015 -3410 1035
rect -3390 1015 -3320 1035
rect -3300 1015 -3230 1035
rect -3210 1015 -3140 1035
rect -3120 1015 -3050 1035
rect -3030 1015 -2960 1035
rect -2940 1015 -2870 1035
rect -2850 1015 -2780 1035
rect -2760 1015 -2690 1035
rect -2670 1015 -2600 1035
rect -2580 1015 -2510 1035
rect -2490 1015 -2420 1035
rect -2400 1015 -2330 1035
rect -2310 1015 -2240 1035
rect -2220 1015 -2150 1035
rect -2130 1015 -2060 1035
rect -2040 1015 -1970 1035
rect -1950 1015 -1880 1035
rect -1860 1015 -1790 1035
rect -1770 1015 -1700 1035
rect -1680 1015 -1610 1035
rect -1590 1015 -1520 1035
rect -1500 1015 -1430 1035
rect -1410 1015 -1340 1035
rect -1320 1015 -1250 1035
rect -1230 1015 -1160 1035
rect -1140 1015 -1070 1035
rect -1050 1015 -980 1035
rect -960 1015 -890 1035
rect -870 1015 -800 1035
rect -780 1015 -710 1035
rect -690 1015 -620 1035
rect -600 1015 -530 1035
rect -510 1015 -440 1035
rect -420 1015 -350 1035
rect -330 1015 -260 1035
rect -240 1015 -170 1035
rect -150 1015 -80 1035
rect -60 1015 45 1035
rect -11615 960 -11510 980
rect -11490 960 -11420 980
rect -11400 960 -11330 980
rect -11310 960 -11240 980
rect -11220 960 -11150 980
rect -11130 960 -11060 980
rect -11040 960 -10970 980
rect -10950 960 -10880 980
rect -10860 960 -10790 980
rect -10770 960 -10700 980
rect -10680 960 -10610 980
rect -10590 960 -10520 980
rect -10500 960 -10430 980
rect -10410 960 -10340 980
rect -10320 960 -10250 980
rect -10230 960 -10160 980
rect -10140 960 -10070 980
rect -10050 960 -9980 980
rect -9960 960 -9890 980
rect -9870 960 -9800 980
rect -9780 960 -9710 980
rect -9690 960 -9620 980
rect -9600 960 -9530 980
rect -9510 960 -9440 980
rect -9420 960 -9350 980
rect -9330 960 -9260 980
rect -9240 960 -9170 980
rect -9150 960 -9080 980
rect -9060 960 -8990 980
rect -8970 960 -8900 980
rect -8880 960 -8810 980
rect -8790 960 -8720 980
rect -8700 960 -8630 980
rect -8610 960 -8540 980
rect -8520 960 -8450 980
rect -8430 960 -8360 980
rect -8340 960 -8270 980
rect -8250 960 -8180 980
rect -8160 960 -8090 980
rect -8070 960 -8000 980
rect -7980 960 -7910 980
rect -7890 960 -7820 980
rect -7800 960 -7730 980
rect -7710 960 -7640 980
rect -7620 960 -7550 980
rect -7530 960 -7460 980
rect -7440 960 -7370 980
rect -7350 960 -7280 980
rect -7260 960 -7190 980
rect -7170 960 -7100 980
rect -7080 960 -7010 980
rect -6990 960 -6920 980
rect -6900 960 -6830 980
rect -6810 960 -6740 980
rect -6720 960 -6650 980
rect -6630 960 -6560 980
rect -6540 960 -6470 980
rect -6450 960 -6380 980
rect -6360 960 -6290 980
rect -6270 960 -6200 980
rect -6180 960 -6110 980
rect -6090 960 -6020 980
rect -6000 960 -5930 980
rect -5910 960 -5840 980
rect -5820 960 -5750 980
rect -5730 960 -5660 980
rect -5640 960 -5570 980
rect -5550 960 -5480 980
rect -5460 960 -5390 980
rect -5370 960 -5300 980
rect -5280 960 -5210 980
rect -5190 960 -5120 980
rect -5100 960 -5030 980
rect -5010 960 -4940 980
rect -4920 960 -4850 980
rect -4830 960 -4760 980
rect -4740 960 -4670 980
rect -4650 960 -4580 980
rect -4560 960 -4490 980
rect -4470 960 -4400 980
rect -4380 960 -4310 980
rect -4290 960 -4220 980
rect -4200 960 -4130 980
rect -4110 960 -4040 980
rect -4020 960 -3950 980
rect -3930 960 -3860 980
rect -3840 960 -3770 980
rect -3750 960 -3680 980
rect -3660 960 -3590 980
rect -3570 960 -3500 980
rect -3480 960 -3410 980
rect -3390 960 -3320 980
rect -3300 960 -3230 980
rect -3210 960 -3140 980
rect -3120 960 -3050 980
rect -3030 960 -2960 980
rect -2940 960 -2870 980
rect -2850 960 -2780 980
rect -2760 960 -2690 980
rect -2670 960 -2600 980
rect -2580 960 -2510 980
rect -2490 960 -2420 980
rect -2400 960 -2330 980
rect -2310 960 -2240 980
rect -2220 960 -2150 980
rect -2130 960 -2060 980
rect -2040 960 -1970 980
rect -1950 960 -1880 980
rect -1860 960 -1790 980
rect -1770 960 -1700 980
rect -1680 960 -1610 980
rect -1590 960 -1520 980
rect -1500 960 -1430 980
rect -1410 960 -1340 980
rect -1320 960 -1250 980
rect -1230 960 -1160 980
rect -1140 960 -1070 980
rect -1050 960 -980 980
rect -960 960 -890 980
rect -870 960 -800 980
rect -780 960 -710 980
rect -690 960 -620 980
rect -600 960 -530 980
rect -510 960 -440 980
rect -420 960 -350 980
rect -330 960 -260 980
rect -240 960 -170 980
rect -150 960 -80 980
rect -60 960 45 980
rect -11615 760 -11595 960
rect 25 760 45 960
rect -11615 740 -11510 760
rect -11490 740 -11420 760
rect -11400 740 -11330 760
rect -11310 740 -11240 760
rect -11220 740 -11150 760
rect -11130 740 -11060 760
rect -11040 740 -10970 760
rect -10950 740 -10880 760
rect -10860 740 -10790 760
rect -10770 740 -10700 760
rect -10680 740 -10610 760
rect -10590 740 -10520 760
rect -10500 740 -10430 760
rect -10410 740 -10340 760
rect -10320 740 -10250 760
rect -10230 740 -10160 760
rect -10140 740 -10070 760
rect -10050 740 -9980 760
rect -9960 740 -9890 760
rect -9870 740 -9800 760
rect -9780 740 -9710 760
rect -9690 740 -9620 760
rect -9600 740 -9530 760
rect -9510 740 -9440 760
rect -9420 740 -9350 760
rect -9330 740 -9260 760
rect -9240 740 -9170 760
rect -9150 740 -9080 760
rect -9060 740 -8990 760
rect -8970 740 -8900 760
rect -8880 740 -8810 760
rect -8790 740 -8720 760
rect -8700 740 -8630 760
rect -8610 740 -8540 760
rect -8520 740 -8450 760
rect -8430 740 -8360 760
rect -8340 740 -8270 760
rect -8250 740 -8180 760
rect -8160 740 -8090 760
rect -8070 740 -8000 760
rect -7980 740 -7910 760
rect -7890 740 -7820 760
rect -7800 740 -7730 760
rect -7710 740 -7640 760
rect -7620 740 -7550 760
rect -7530 740 -7460 760
rect -7440 740 -7370 760
rect -7350 740 -7280 760
rect -7260 740 -7190 760
rect -7170 740 -7100 760
rect -7080 740 -7010 760
rect -6990 740 -6920 760
rect -6900 740 -6830 760
rect -6810 740 -6740 760
rect -6720 740 -6650 760
rect -6630 740 -6560 760
rect -6540 740 -6470 760
rect -6450 740 -6380 760
rect -6360 740 -6290 760
rect -6270 740 -6200 760
rect -6180 740 -6110 760
rect -6090 740 -6020 760
rect -6000 740 -5930 760
rect -5910 740 -5840 760
rect -5820 740 -5750 760
rect -5730 740 -5660 760
rect -5640 740 -5570 760
rect -5550 740 -5480 760
rect -5460 740 -5390 760
rect -5370 740 -5300 760
rect -5280 740 -5210 760
rect -5190 740 -5120 760
rect -5100 740 -5030 760
rect -5010 740 -4940 760
rect -4920 740 -4850 760
rect -4830 740 -4760 760
rect -4740 740 -4670 760
rect -4650 740 -4580 760
rect -4560 740 -4490 760
rect -4470 740 -4400 760
rect -4380 740 -4310 760
rect -4290 740 -4220 760
rect -4200 740 -4130 760
rect -4110 740 -4040 760
rect -4020 740 -3950 760
rect -3930 740 -3860 760
rect -3840 740 -3770 760
rect -3750 740 -3680 760
rect -3660 740 -3590 760
rect -3570 740 -3500 760
rect -3480 740 -3410 760
rect -3390 740 -3320 760
rect -3300 740 -3230 760
rect -3210 740 -3140 760
rect -3120 740 -3050 760
rect -3030 740 -2960 760
rect -2940 740 -2870 760
rect -2850 740 -2780 760
rect -2760 740 -2690 760
rect -2670 740 -2600 760
rect -2580 740 -2510 760
rect -2490 740 -2420 760
rect -2400 740 -2330 760
rect -2310 740 -2240 760
rect -2220 740 -2150 760
rect -2130 740 -2060 760
rect -2040 740 -1970 760
rect -1950 740 -1880 760
rect -1860 740 -1790 760
rect -1770 740 -1700 760
rect -1680 740 -1610 760
rect -1590 740 -1520 760
rect -1500 740 -1430 760
rect -1410 740 -1340 760
rect -1320 740 -1250 760
rect -1230 740 -1160 760
rect -1140 740 -1070 760
rect -1050 740 -980 760
rect -960 740 -890 760
rect -870 740 -800 760
rect -780 740 -710 760
rect -690 740 -620 760
rect -600 740 -530 760
rect -510 740 -440 760
rect -420 740 -350 760
rect -330 740 -260 760
rect -240 740 -170 760
rect -150 740 -80 760
rect -60 740 45 760
<< psubdiffcont >>
rect -11510 1975 -11490 1995
rect -11420 1975 -11400 1995
rect -11330 1975 -11310 1995
rect -11240 1975 -11220 1995
rect -11150 1975 -11130 1995
rect -11060 1975 -11040 1995
rect -10970 1975 -10950 1995
rect -10880 1975 -10860 1995
rect -10790 1975 -10770 1995
rect -10700 1975 -10680 1995
rect -10610 1975 -10590 1995
rect -10520 1975 -10500 1995
rect -10430 1975 -10410 1995
rect -10340 1975 -10320 1995
rect -10250 1975 -10230 1995
rect -10160 1975 -10140 1995
rect -10070 1975 -10050 1995
rect -9980 1975 -9960 1995
rect -9890 1975 -9870 1995
rect -9800 1975 -9780 1995
rect -9710 1975 -9690 1995
rect -9620 1975 -9600 1995
rect -9530 1975 -9510 1995
rect -9440 1975 -9420 1995
rect -9350 1975 -9330 1995
rect -9260 1975 -9240 1995
rect -9170 1975 -9150 1995
rect -9080 1975 -9060 1995
rect -8990 1975 -8970 1995
rect -8900 1975 -8880 1995
rect -8810 1975 -8790 1995
rect -8720 1975 -8700 1995
rect -8630 1975 -8610 1995
rect -8540 1975 -8520 1995
rect -8450 1975 -8430 1995
rect -8360 1975 -8340 1995
rect -8270 1975 -8250 1995
rect -8180 1975 -8160 1995
rect -8090 1975 -8070 1995
rect -8000 1975 -7980 1995
rect -7910 1975 -7890 1995
rect -7820 1975 -7800 1995
rect -7730 1975 -7710 1995
rect -7640 1975 -7620 1995
rect -7550 1975 -7530 1995
rect -7460 1975 -7440 1995
rect -7370 1975 -7350 1995
rect -7280 1975 -7260 1995
rect -7190 1975 -7170 1995
rect -7100 1975 -7080 1995
rect -7010 1975 -6990 1995
rect -6920 1975 -6900 1995
rect -6830 1975 -6810 1995
rect -6740 1975 -6720 1995
rect -6650 1975 -6630 1995
rect -6560 1975 -6540 1995
rect -6470 1975 -6450 1995
rect -6380 1975 -6360 1995
rect -6290 1975 -6270 1995
rect -6200 1975 -6180 1995
rect -6110 1975 -6090 1995
rect -6020 1975 -6000 1995
rect -5930 1975 -5910 1995
rect -5840 1975 -5820 1995
rect -5750 1975 -5730 1995
rect -5660 1975 -5640 1995
rect -5570 1975 -5550 1995
rect -5480 1975 -5460 1995
rect -5390 1975 -5370 1995
rect -5300 1975 -5280 1995
rect -5210 1975 -5190 1995
rect -5120 1975 -5100 1995
rect -5030 1975 -5010 1995
rect -4940 1975 -4920 1995
rect -4850 1975 -4830 1995
rect -4760 1975 -4740 1995
rect -4670 1975 -4650 1995
rect -4580 1975 -4560 1995
rect -4490 1975 -4470 1995
rect -4400 1975 -4380 1995
rect -4310 1975 -4290 1995
rect -4220 1975 -4200 1995
rect -4130 1975 -4110 1995
rect -4040 1975 -4020 1995
rect -3950 1975 -3930 1995
rect -3860 1975 -3840 1995
rect -3770 1975 -3750 1995
rect -3680 1975 -3660 1995
rect -3590 1975 -3570 1995
rect -3500 1975 -3480 1995
rect -3410 1975 -3390 1995
rect -3320 1975 -3300 1995
rect -3230 1975 -3210 1995
rect -3140 1975 -3120 1995
rect -3050 1975 -3030 1995
rect -2960 1975 -2940 1995
rect -2870 1975 -2850 1995
rect -2780 1975 -2760 1995
rect -2690 1975 -2670 1995
rect -2600 1975 -2580 1995
rect -2510 1975 -2490 1995
rect -2420 1975 -2400 1995
rect -2330 1975 -2310 1995
rect -2240 1975 -2220 1995
rect -2150 1975 -2130 1995
rect -2060 1975 -2040 1995
rect -1970 1975 -1950 1995
rect -1880 1975 -1860 1995
rect -1790 1975 -1770 1995
rect -1700 1975 -1680 1995
rect -1610 1975 -1590 1995
rect -1520 1975 -1500 1995
rect -1430 1975 -1410 1995
rect -1340 1975 -1320 1995
rect -1250 1975 -1230 1995
rect -1160 1975 -1140 1995
rect -1070 1975 -1050 1995
rect -980 1975 -960 1995
rect -890 1975 -870 1995
rect -800 1975 -780 1995
rect -710 1975 -690 1995
rect -620 1975 -600 1995
rect -530 1975 -510 1995
rect -440 1975 -420 1995
rect -350 1975 -330 1995
rect -260 1975 -240 1995
rect -170 1975 -150 1995
rect -80 1975 -60 1995
rect -11510 1755 -11490 1775
rect -11420 1755 -11400 1775
rect -11330 1755 -11310 1775
rect -11240 1755 -11220 1775
rect -11150 1755 -11130 1775
rect -11060 1755 -11040 1775
rect -10970 1755 -10950 1775
rect -10880 1755 -10860 1775
rect -10790 1755 -10770 1775
rect -10700 1755 -10680 1775
rect -10610 1755 -10590 1775
rect -10520 1755 -10500 1775
rect -10430 1755 -10410 1775
rect -10340 1755 -10320 1775
rect -10250 1755 -10230 1775
rect -10160 1755 -10140 1775
rect -10070 1755 -10050 1775
rect -9980 1755 -9960 1775
rect -9890 1755 -9870 1775
rect -9800 1755 -9780 1775
rect -9710 1755 -9690 1775
rect -9620 1755 -9600 1775
rect -9530 1755 -9510 1775
rect -9440 1755 -9420 1775
rect -9350 1755 -9330 1775
rect -9260 1755 -9240 1775
rect -9170 1755 -9150 1775
rect -9080 1755 -9060 1775
rect -8990 1755 -8970 1775
rect -8900 1755 -8880 1775
rect -8810 1755 -8790 1775
rect -8720 1755 -8700 1775
rect -8630 1755 -8610 1775
rect -8540 1755 -8520 1775
rect -8450 1755 -8430 1775
rect -8360 1755 -8340 1775
rect -8270 1755 -8250 1775
rect -8180 1755 -8160 1775
rect -8090 1755 -8070 1775
rect -8000 1755 -7980 1775
rect -7910 1755 -7890 1775
rect -7820 1755 -7800 1775
rect -7730 1755 -7710 1775
rect -7640 1755 -7620 1775
rect -7550 1755 -7530 1775
rect -7460 1755 -7440 1775
rect -7370 1755 -7350 1775
rect -7280 1755 -7260 1775
rect -7190 1755 -7170 1775
rect -7100 1755 -7080 1775
rect -7010 1755 -6990 1775
rect -6920 1755 -6900 1775
rect -6830 1755 -6810 1775
rect -6740 1755 -6720 1775
rect -6650 1755 -6630 1775
rect -6560 1755 -6540 1775
rect -6470 1755 -6450 1775
rect -6380 1755 -6360 1775
rect -6290 1755 -6270 1775
rect -6200 1755 -6180 1775
rect -6110 1755 -6090 1775
rect -6020 1755 -6000 1775
rect -5930 1755 -5910 1775
rect -5840 1755 -5820 1775
rect -5750 1755 -5730 1775
rect -5660 1755 -5640 1775
rect -5570 1755 -5550 1775
rect -5480 1755 -5460 1775
rect -5390 1755 -5370 1775
rect -5300 1755 -5280 1775
rect -5210 1755 -5190 1775
rect -5120 1755 -5100 1775
rect -5030 1755 -5010 1775
rect -4940 1755 -4920 1775
rect -4850 1755 -4830 1775
rect -4760 1755 -4740 1775
rect -4670 1755 -4650 1775
rect -4580 1755 -4560 1775
rect -4490 1755 -4470 1775
rect -4400 1755 -4380 1775
rect -4310 1755 -4290 1775
rect -4220 1755 -4200 1775
rect -4130 1755 -4110 1775
rect -4040 1755 -4020 1775
rect -3950 1755 -3930 1775
rect -3860 1755 -3840 1775
rect -3770 1755 -3750 1775
rect -3680 1755 -3660 1775
rect -3590 1755 -3570 1775
rect -3500 1755 -3480 1775
rect -3410 1755 -3390 1775
rect -3320 1755 -3300 1775
rect -3230 1755 -3210 1775
rect -3140 1755 -3120 1775
rect -3050 1755 -3030 1775
rect -2960 1755 -2940 1775
rect -2870 1755 -2850 1775
rect -2780 1755 -2760 1775
rect -2690 1755 -2670 1775
rect -2600 1755 -2580 1775
rect -2510 1755 -2490 1775
rect -2420 1755 -2400 1775
rect -2330 1755 -2310 1775
rect -2240 1755 -2220 1775
rect -2150 1755 -2130 1775
rect -2060 1755 -2040 1775
rect -1970 1755 -1950 1775
rect -1880 1755 -1860 1775
rect -1790 1755 -1770 1775
rect -1700 1755 -1680 1775
rect -1610 1755 -1590 1775
rect -1520 1755 -1500 1775
rect -1430 1755 -1410 1775
rect -1340 1755 -1320 1775
rect -1250 1755 -1230 1775
rect -1160 1755 -1140 1775
rect -1070 1755 -1050 1775
rect -980 1755 -960 1775
rect -890 1755 -870 1775
rect -800 1755 -780 1775
rect -710 1755 -690 1775
rect -620 1755 -600 1775
rect -530 1755 -510 1775
rect -440 1755 -420 1775
rect -350 1755 -330 1775
rect -260 1755 -240 1775
rect -170 1755 -150 1775
rect -80 1755 -60 1775
rect -11510 1315 -11490 1335
rect -11420 1315 -11400 1335
rect -11330 1315 -11310 1335
rect -11240 1315 -11220 1335
rect -11150 1315 -11130 1335
rect -11060 1315 -11040 1335
rect -10970 1315 -10950 1335
rect -10880 1315 -10860 1335
rect -10790 1315 -10770 1335
rect -10700 1315 -10680 1335
rect -10610 1315 -10590 1335
rect -10520 1315 -10500 1335
rect -10430 1315 -10410 1335
rect -10340 1315 -10320 1335
rect -10250 1315 -10230 1335
rect -10160 1315 -10140 1335
rect -10070 1315 -10050 1335
rect -9980 1315 -9960 1335
rect -9890 1315 -9870 1335
rect -9800 1315 -9780 1335
rect -9710 1315 -9690 1335
rect -9620 1315 -9600 1335
rect -9530 1315 -9510 1335
rect -9440 1315 -9420 1335
rect -9350 1315 -9330 1335
rect -9260 1315 -9240 1335
rect -9170 1315 -9150 1335
rect -9080 1315 -9060 1335
rect -8990 1315 -8970 1335
rect -8900 1315 -8880 1335
rect -8810 1315 -8790 1335
rect -8720 1315 -8700 1335
rect -8630 1315 -8610 1335
rect -8540 1315 -8520 1335
rect -8450 1315 -8430 1335
rect -8360 1315 -8340 1335
rect -8270 1315 -8250 1335
rect -8180 1315 -8160 1335
rect -8090 1315 -8070 1335
rect -8000 1315 -7980 1335
rect -7910 1315 -7890 1335
rect -7820 1315 -7800 1335
rect -7730 1315 -7710 1335
rect -7640 1315 -7620 1335
rect -7550 1315 -7530 1335
rect -7460 1315 -7440 1335
rect -7370 1315 -7350 1335
rect -7280 1315 -7260 1335
rect -7190 1315 -7170 1335
rect -7100 1315 -7080 1335
rect -7010 1315 -6990 1335
rect -6920 1315 -6900 1335
rect -6830 1315 -6810 1335
rect -6740 1315 -6720 1335
rect -6650 1315 -6630 1335
rect -6560 1315 -6540 1335
rect -6470 1315 -6450 1335
rect -6380 1315 -6360 1335
rect -6290 1315 -6270 1335
rect -6200 1315 -6180 1335
rect -6110 1315 -6090 1335
rect -6020 1315 -6000 1335
rect -5930 1315 -5910 1335
rect -5840 1315 -5820 1335
rect -5750 1315 -5730 1335
rect -5660 1315 -5640 1335
rect -5570 1315 -5550 1335
rect -5480 1315 -5460 1335
rect -5390 1315 -5370 1335
rect -5300 1315 -5280 1335
rect -5210 1315 -5190 1335
rect -5120 1315 -5100 1335
rect -5030 1315 -5010 1335
rect -4940 1315 -4920 1335
rect -4850 1315 -4830 1335
rect -4760 1315 -4740 1335
rect -4670 1315 -4650 1335
rect -4580 1315 -4560 1335
rect -4490 1315 -4470 1335
rect -4400 1315 -4380 1335
rect -4310 1315 -4290 1335
rect -4220 1315 -4200 1335
rect -4130 1315 -4110 1335
rect -4040 1315 -4020 1335
rect -3950 1315 -3930 1335
rect -3860 1315 -3840 1335
rect -3770 1315 -3750 1335
rect -3680 1315 -3660 1335
rect -3590 1315 -3570 1335
rect -3500 1315 -3480 1335
rect -3410 1315 -3390 1335
rect -3320 1315 -3300 1335
rect -3230 1315 -3210 1335
rect -3140 1315 -3120 1335
rect -3050 1315 -3030 1335
rect -2960 1315 -2940 1335
rect -2870 1315 -2850 1335
rect -2780 1315 -2760 1335
rect -2690 1315 -2670 1335
rect -2600 1315 -2580 1335
rect -2510 1315 -2490 1335
rect -2420 1315 -2400 1335
rect -2330 1315 -2310 1335
rect -2240 1315 -2220 1335
rect -2150 1315 -2130 1335
rect -2060 1315 -2040 1335
rect -1970 1315 -1950 1335
rect -1880 1315 -1860 1335
rect -1790 1315 -1770 1335
rect -1700 1315 -1680 1335
rect -1610 1315 -1590 1335
rect -1520 1315 -1500 1335
rect -1430 1315 -1410 1335
rect -1340 1315 -1320 1335
rect -1250 1315 -1230 1335
rect -1160 1315 -1140 1335
rect -1070 1315 -1050 1335
rect -980 1315 -960 1335
rect -890 1315 -870 1335
rect -800 1315 -780 1335
rect -710 1315 -690 1335
rect -620 1315 -600 1335
rect -530 1315 -510 1335
rect -440 1315 -420 1335
rect -350 1315 -330 1335
rect -260 1315 -240 1335
rect -170 1315 -150 1335
rect -80 1315 -60 1335
rect -11510 660 -11490 680
rect -11420 660 -11400 680
rect -11330 660 -11310 680
rect -11240 660 -11220 680
rect -11150 660 -11130 680
rect -11060 660 -11040 680
rect -10970 660 -10950 680
rect -10880 660 -10860 680
rect -10790 660 -10770 680
rect -10700 660 -10680 680
rect -10610 660 -10590 680
rect -10520 660 -10500 680
rect -10430 660 -10410 680
rect -10340 660 -10320 680
rect -10250 660 -10230 680
rect -10160 660 -10140 680
rect -10070 660 -10050 680
rect -9980 660 -9960 680
rect -9890 660 -9870 680
rect -9800 660 -9780 680
rect -9710 660 -9690 680
rect -9620 660 -9600 680
rect -9530 660 -9510 680
rect -9440 660 -9420 680
rect -9350 660 -9330 680
rect -9260 660 -9240 680
rect -9170 660 -9150 680
rect -9080 660 -9060 680
rect -8990 660 -8970 680
rect -8900 660 -8880 680
rect -8810 660 -8790 680
rect -8720 660 -8700 680
rect -8630 660 -8610 680
rect -8540 660 -8520 680
rect -8450 660 -8430 680
rect -8360 660 -8340 680
rect -8270 660 -8250 680
rect -8180 660 -8160 680
rect -8090 660 -8070 680
rect -8000 660 -7980 680
rect -7910 660 -7890 680
rect -7820 660 -7800 680
rect -7730 660 -7710 680
rect -7640 660 -7620 680
rect -7550 660 -7530 680
rect -7460 660 -7440 680
rect -7370 660 -7350 680
rect -7280 660 -7260 680
rect -7190 660 -7170 680
rect -7100 660 -7080 680
rect -7010 660 -6990 680
rect -6920 660 -6900 680
rect -6830 660 -6810 680
rect -6740 660 -6720 680
rect -6650 660 -6630 680
rect -6560 660 -6540 680
rect -6470 660 -6450 680
rect -6380 660 -6360 680
rect -6290 660 -6270 680
rect -6200 660 -6180 680
rect -6110 660 -6090 680
rect -6020 660 -6000 680
rect -5930 660 -5910 680
rect -5840 660 -5820 680
rect -5750 660 -5730 680
rect -5660 660 -5640 680
rect -5570 660 -5550 680
rect -5480 660 -5460 680
rect -5390 660 -5370 680
rect -5300 660 -5280 680
rect -5210 660 -5190 680
rect -5120 660 -5100 680
rect -5030 660 -5010 680
rect -4940 660 -4920 680
rect -4850 660 -4830 680
rect -4760 660 -4740 680
rect -4670 660 -4650 680
rect -4580 660 -4560 680
rect -4490 660 -4470 680
rect -4400 660 -4380 680
rect -4310 660 -4290 680
rect -4220 660 -4200 680
rect -4130 660 -4110 680
rect -4040 660 -4020 680
rect -3950 660 -3930 680
rect -3860 660 -3840 680
rect -3770 660 -3750 680
rect -3680 660 -3660 680
rect -3590 660 -3570 680
rect -3500 660 -3480 680
rect -3410 660 -3390 680
rect -3320 660 -3300 680
rect -3230 660 -3210 680
rect -3140 660 -3120 680
rect -3050 660 -3030 680
rect -2960 660 -2940 680
rect -2870 660 -2850 680
rect -2780 660 -2760 680
rect -2690 660 -2670 680
rect -2600 660 -2580 680
rect -2510 660 -2490 680
rect -2420 660 -2400 680
rect -2330 660 -2310 680
rect -2240 660 -2220 680
rect -2150 660 -2130 680
rect -2060 660 -2040 680
rect -1970 660 -1950 680
rect -1880 660 -1860 680
rect -1790 660 -1770 680
rect -1700 660 -1680 680
rect -1610 660 -1590 680
rect -1520 660 -1500 680
rect -1430 660 -1410 680
rect -1340 660 -1320 680
rect -1250 660 -1230 680
rect -1160 660 -1140 680
rect -1070 660 -1050 680
rect -980 660 -960 680
rect -890 660 -870 680
rect -800 660 -780 680
rect -710 660 -690 680
rect -620 660 -600 680
rect -530 660 -510 680
rect -440 660 -420 680
rect -350 660 -330 680
rect -260 660 -240 680
rect -170 660 -150 680
rect -80 660 -60 680
rect -11510 220 -11490 240
rect -11420 220 -11400 240
rect -11330 220 -11310 240
rect -11240 220 -11220 240
rect -11150 220 -11130 240
rect -11060 220 -11040 240
rect -10970 220 -10950 240
rect -10880 220 -10860 240
rect -10790 220 -10770 240
rect -10700 220 -10680 240
rect -10610 220 -10590 240
rect -10520 220 -10500 240
rect -10430 220 -10410 240
rect -10340 220 -10320 240
rect -10250 220 -10230 240
rect -10160 220 -10140 240
rect -10070 220 -10050 240
rect -9980 220 -9960 240
rect -9890 220 -9870 240
rect -9800 220 -9780 240
rect -9710 220 -9690 240
rect -9620 220 -9600 240
rect -9530 220 -9510 240
rect -9440 220 -9420 240
rect -9350 220 -9330 240
rect -9260 220 -9240 240
rect -9170 220 -9150 240
rect -9080 220 -9060 240
rect -8990 220 -8970 240
rect -8900 220 -8880 240
rect -8810 220 -8790 240
rect -8720 220 -8700 240
rect -8630 220 -8610 240
rect -8540 220 -8520 240
rect -8450 220 -8430 240
rect -8360 220 -8340 240
rect -8270 220 -8250 240
rect -8180 220 -8160 240
rect -8090 220 -8070 240
rect -8000 220 -7980 240
rect -7910 220 -7890 240
rect -7820 220 -7800 240
rect -7730 220 -7710 240
rect -7640 220 -7620 240
rect -7550 220 -7530 240
rect -7460 220 -7440 240
rect -7370 220 -7350 240
rect -7280 220 -7260 240
rect -7190 220 -7170 240
rect -7100 220 -7080 240
rect -7010 220 -6990 240
rect -6920 220 -6900 240
rect -6830 220 -6810 240
rect -6740 220 -6720 240
rect -6650 220 -6630 240
rect -6560 220 -6540 240
rect -6470 220 -6450 240
rect -6380 220 -6360 240
rect -6290 220 -6270 240
rect -6200 220 -6180 240
rect -6110 220 -6090 240
rect -6020 220 -6000 240
rect -5930 220 -5910 240
rect -5840 220 -5820 240
rect -5750 220 -5730 240
rect -5660 220 -5640 240
rect -5570 220 -5550 240
rect -5480 220 -5460 240
rect -5390 220 -5370 240
rect -5300 220 -5280 240
rect -5210 220 -5190 240
rect -5120 220 -5100 240
rect -5030 220 -5010 240
rect -4940 220 -4920 240
rect -4850 220 -4830 240
rect -4760 220 -4740 240
rect -4670 220 -4650 240
rect -4580 220 -4560 240
rect -4490 220 -4470 240
rect -4400 220 -4380 240
rect -4310 220 -4290 240
rect -4220 220 -4200 240
rect -4130 220 -4110 240
rect -4040 220 -4020 240
rect -3950 220 -3930 240
rect -3860 220 -3840 240
rect -3770 220 -3750 240
rect -3680 220 -3660 240
rect -3590 220 -3570 240
rect -3500 220 -3480 240
rect -3410 220 -3390 240
rect -3320 220 -3300 240
rect -3230 220 -3210 240
rect -3140 220 -3120 240
rect -3050 220 -3030 240
rect -2960 220 -2940 240
rect -2870 220 -2850 240
rect -2780 220 -2760 240
rect -2690 220 -2670 240
rect -2600 220 -2580 240
rect -2510 220 -2490 240
rect -2420 220 -2400 240
rect -2330 220 -2310 240
rect -2240 220 -2220 240
rect -2150 220 -2130 240
rect -2060 220 -2040 240
rect -1970 220 -1950 240
rect -1880 220 -1860 240
rect -1790 220 -1770 240
rect -1700 220 -1680 240
rect -1610 220 -1590 240
rect -1520 220 -1500 240
rect -1430 220 -1410 240
rect -1340 220 -1320 240
rect -1250 220 -1230 240
rect -1160 220 -1140 240
rect -1070 220 -1050 240
rect -980 220 -960 240
rect -890 220 -870 240
rect -800 220 -780 240
rect -710 220 -690 240
rect -620 220 -600 240
rect -530 220 -510 240
rect -440 220 -420 240
rect -350 220 -330 240
rect -260 220 -240 240
rect -170 220 -150 240
rect -80 220 -60 240
rect -11510 0 -11490 20
rect -11420 0 -11400 20
rect -11330 0 -11310 20
rect -11240 0 -11220 20
rect -11150 0 -11130 20
rect -11060 0 -11040 20
rect -10970 0 -10950 20
rect -10880 0 -10860 20
rect -10790 0 -10770 20
rect -10700 0 -10680 20
rect -10610 0 -10590 20
rect -10520 0 -10500 20
rect -10430 0 -10410 20
rect -10340 0 -10320 20
rect -10250 0 -10230 20
rect -10160 0 -10140 20
rect -10070 0 -10050 20
rect -9980 0 -9960 20
rect -9890 0 -9870 20
rect -9800 0 -9780 20
rect -9710 0 -9690 20
rect -9620 0 -9600 20
rect -9530 0 -9510 20
rect -9440 0 -9420 20
rect -9350 0 -9330 20
rect -9260 0 -9240 20
rect -9170 0 -9150 20
rect -9080 0 -9060 20
rect -8990 0 -8970 20
rect -8900 0 -8880 20
rect -8810 0 -8790 20
rect -8720 0 -8700 20
rect -8630 0 -8610 20
rect -8540 0 -8520 20
rect -8450 0 -8430 20
rect -8360 0 -8340 20
rect -8270 0 -8250 20
rect -8180 0 -8160 20
rect -8090 0 -8070 20
rect -8000 0 -7980 20
rect -7910 0 -7890 20
rect -7820 0 -7800 20
rect -7730 0 -7710 20
rect -7640 0 -7620 20
rect -7550 0 -7530 20
rect -7460 0 -7440 20
rect -7370 0 -7350 20
rect -7280 0 -7260 20
rect -7190 0 -7170 20
rect -7100 0 -7080 20
rect -7010 0 -6990 20
rect -6920 0 -6900 20
rect -6830 0 -6810 20
rect -6740 0 -6720 20
rect -6650 0 -6630 20
rect -6560 0 -6540 20
rect -6470 0 -6450 20
rect -6380 0 -6360 20
rect -6290 0 -6270 20
rect -6200 0 -6180 20
rect -6110 0 -6090 20
rect -6020 0 -6000 20
rect -5930 0 -5910 20
rect -5840 0 -5820 20
rect -5750 0 -5730 20
rect -5660 0 -5640 20
rect -5570 0 -5550 20
rect -5480 0 -5460 20
rect -5390 0 -5370 20
rect -5300 0 -5280 20
rect -5210 0 -5190 20
rect -5120 0 -5100 20
rect -5030 0 -5010 20
rect -4940 0 -4920 20
rect -4850 0 -4830 20
rect -4760 0 -4740 20
rect -4670 0 -4650 20
rect -4580 0 -4560 20
rect -4490 0 -4470 20
rect -4400 0 -4380 20
rect -4310 0 -4290 20
rect -4220 0 -4200 20
rect -4130 0 -4110 20
rect -4040 0 -4020 20
rect -3950 0 -3930 20
rect -3860 0 -3840 20
rect -3770 0 -3750 20
rect -3680 0 -3660 20
rect -3590 0 -3570 20
rect -3500 0 -3480 20
rect -3410 0 -3390 20
rect -3320 0 -3300 20
rect -3230 0 -3210 20
rect -3140 0 -3120 20
rect -3050 0 -3030 20
rect -2960 0 -2940 20
rect -2870 0 -2850 20
rect -2780 0 -2760 20
rect -2690 0 -2670 20
rect -2600 0 -2580 20
rect -2510 0 -2490 20
rect -2420 0 -2400 20
rect -2330 0 -2310 20
rect -2240 0 -2220 20
rect -2150 0 -2130 20
rect -2060 0 -2040 20
rect -1970 0 -1950 20
rect -1880 0 -1860 20
rect -1790 0 -1770 20
rect -1700 0 -1680 20
rect -1610 0 -1590 20
rect -1520 0 -1500 20
rect -1430 0 -1410 20
rect -1340 0 -1320 20
rect -1250 0 -1230 20
rect -1160 0 -1140 20
rect -1070 0 -1050 20
rect -980 0 -960 20
rect -890 0 -870 20
rect -800 0 -780 20
rect -710 0 -690 20
rect -620 0 -600 20
rect -530 0 -510 20
rect -440 0 -420 20
rect -350 0 -330 20
rect -260 0 -240 20
rect -170 0 -150 20
rect -80 0 -60 20
<< nsubdiffcont >>
rect -11510 1235 -11490 1255
rect -11420 1235 -11400 1255
rect -11330 1235 -11310 1255
rect -11240 1235 -11220 1255
rect -11150 1235 -11130 1255
rect -11060 1235 -11040 1255
rect -10970 1235 -10950 1255
rect -10880 1235 -10860 1255
rect -10790 1235 -10770 1255
rect -10700 1235 -10680 1255
rect -10610 1235 -10590 1255
rect -10520 1235 -10500 1255
rect -10430 1235 -10410 1255
rect -10340 1235 -10320 1255
rect -10250 1235 -10230 1255
rect -10160 1235 -10140 1255
rect -10070 1235 -10050 1255
rect -9980 1235 -9960 1255
rect -9890 1235 -9870 1255
rect -9800 1235 -9780 1255
rect -9710 1235 -9690 1255
rect -9620 1235 -9600 1255
rect -9530 1235 -9510 1255
rect -9440 1235 -9420 1255
rect -9350 1235 -9330 1255
rect -9260 1235 -9240 1255
rect -9170 1235 -9150 1255
rect -9080 1235 -9060 1255
rect -8990 1235 -8970 1255
rect -8900 1235 -8880 1255
rect -8810 1235 -8790 1255
rect -8720 1235 -8700 1255
rect -8630 1235 -8610 1255
rect -8540 1235 -8520 1255
rect -8450 1235 -8430 1255
rect -8360 1235 -8340 1255
rect -8270 1235 -8250 1255
rect -8180 1235 -8160 1255
rect -8090 1235 -8070 1255
rect -8000 1235 -7980 1255
rect -7910 1235 -7890 1255
rect -7820 1235 -7800 1255
rect -7730 1235 -7710 1255
rect -7640 1235 -7620 1255
rect -7550 1235 -7530 1255
rect -7460 1235 -7440 1255
rect -7370 1235 -7350 1255
rect -7280 1235 -7260 1255
rect -7190 1235 -7170 1255
rect -7100 1235 -7080 1255
rect -7010 1235 -6990 1255
rect -6920 1235 -6900 1255
rect -6830 1235 -6810 1255
rect -6740 1235 -6720 1255
rect -6650 1235 -6630 1255
rect -6560 1235 -6540 1255
rect -6470 1235 -6450 1255
rect -6380 1235 -6360 1255
rect -6290 1235 -6270 1255
rect -6200 1235 -6180 1255
rect -6110 1235 -6090 1255
rect -6020 1235 -6000 1255
rect -5930 1235 -5910 1255
rect -5840 1235 -5820 1255
rect -5750 1235 -5730 1255
rect -5660 1235 -5640 1255
rect -5570 1235 -5550 1255
rect -5480 1235 -5460 1255
rect -5390 1235 -5370 1255
rect -5300 1235 -5280 1255
rect -5210 1235 -5190 1255
rect -5120 1235 -5100 1255
rect -5030 1235 -5010 1255
rect -4940 1235 -4920 1255
rect -4850 1235 -4830 1255
rect -4760 1235 -4740 1255
rect -4670 1235 -4650 1255
rect -4580 1235 -4560 1255
rect -4490 1235 -4470 1255
rect -4400 1235 -4380 1255
rect -4310 1235 -4290 1255
rect -4220 1235 -4200 1255
rect -4130 1235 -4110 1255
rect -4040 1235 -4020 1255
rect -3950 1235 -3930 1255
rect -3860 1235 -3840 1255
rect -3770 1235 -3750 1255
rect -3680 1235 -3660 1255
rect -3590 1235 -3570 1255
rect -3500 1235 -3480 1255
rect -3410 1235 -3390 1255
rect -3320 1235 -3300 1255
rect -3230 1235 -3210 1255
rect -3140 1235 -3120 1255
rect -3050 1235 -3030 1255
rect -2960 1235 -2940 1255
rect -2870 1235 -2850 1255
rect -2780 1235 -2760 1255
rect -2690 1235 -2670 1255
rect -2600 1235 -2580 1255
rect -2510 1235 -2490 1255
rect -2420 1235 -2400 1255
rect -2330 1235 -2310 1255
rect -2240 1235 -2220 1255
rect -2150 1235 -2130 1255
rect -2060 1235 -2040 1255
rect -1970 1235 -1950 1255
rect -1880 1235 -1860 1255
rect -1790 1235 -1770 1255
rect -1700 1235 -1680 1255
rect -1610 1235 -1590 1255
rect -1520 1235 -1500 1255
rect -1430 1235 -1410 1255
rect -1340 1235 -1320 1255
rect -1250 1235 -1230 1255
rect -1160 1235 -1140 1255
rect -1070 1235 -1050 1255
rect -980 1235 -960 1255
rect -890 1235 -870 1255
rect -800 1235 -780 1255
rect -710 1235 -690 1255
rect -620 1235 -600 1255
rect -530 1235 -510 1255
rect -440 1235 -420 1255
rect -350 1235 -330 1255
rect -260 1235 -240 1255
rect -170 1235 -150 1255
rect -80 1235 -60 1255
rect -11510 1015 -11490 1035
rect -11420 1015 -11400 1035
rect -11330 1015 -11310 1035
rect -11240 1015 -11220 1035
rect -11150 1015 -11130 1035
rect -11060 1015 -11040 1035
rect -10970 1015 -10950 1035
rect -10880 1015 -10860 1035
rect -10790 1015 -10770 1035
rect -10700 1015 -10680 1035
rect -10610 1015 -10590 1035
rect -10520 1015 -10500 1035
rect -10430 1015 -10410 1035
rect -10340 1015 -10320 1035
rect -10250 1015 -10230 1035
rect -10160 1015 -10140 1035
rect -10070 1015 -10050 1035
rect -9980 1015 -9960 1035
rect -9890 1015 -9870 1035
rect -9800 1015 -9780 1035
rect -9710 1015 -9690 1035
rect -9620 1015 -9600 1035
rect -9530 1015 -9510 1035
rect -9440 1015 -9420 1035
rect -9350 1015 -9330 1035
rect -9260 1015 -9240 1035
rect -9170 1015 -9150 1035
rect -9080 1015 -9060 1035
rect -8990 1015 -8970 1035
rect -8900 1015 -8880 1035
rect -8810 1015 -8790 1035
rect -8720 1015 -8700 1035
rect -8630 1015 -8610 1035
rect -8540 1015 -8520 1035
rect -8450 1015 -8430 1035
rect -8360 1015 -8340 1035
rect -8270 1015 -8250 1035
rect -8180 1015 -8160 1035
rect -8090 1015 -8070 1035
rect -8000 1015 -7980 1035
rect -7910 1015 -7890 1035
rect -7820 1015 -7800 1035
rect -7730 1015 -7710 1035
rect -7640 1015 -7620 1035
rect -7550 1015 -7530 1035
rect -7460 1015 -7440 1035
rect -7370 1015 -7350 1035
rect -7280 1015 -7260 1035
rect -7190 1015 -7170 1035
rect -7100 1015 -7080 1035
rect -7010 1015 -6990 1035
rect -6920 1015 -6900 1035
rect -6830 1015 -6810 1035
rect -6740 1015 -6720 1035
rect -6650 1015 -6630 1035
rect -6560 1015 -6540 1035
rect -6470 1015 -6450 1035
rect -6380 1015 -6360 1035
rect -6290 1015 -6270 1035
rect -6200 1015 -6180 1035
rect -6110 1015 -6090 1035
rect -6020 1015 -6000 1035
rect -5930 1015 -5910 1035
rect -5840 1015 -5820 1035
rect -5750 1015 -5730 1035
rect -5660 1015 -5640 1035
rect -5570 1015 -5550 1035
rect -5480 1015 -5460 1035
rect -5390 1015 -5370 1035
rect -5300 1015 -5280 1035
rect -5210 1015 -5190 1035
rect -5120 1015 -5100 1035
rect -5030 1015 -5010 1035
rect -4940 1015 -4920 1035
rect -4850 1015 -4830 1035
rect -4760 1015 -4740 1035
rect -4670 1015 -4650 1035
rect -4580 1015 -4560 1035
rect -4490 1015 -4470 1035
rect -4400 1015 -4380 1035
rect -4310 1015 -4290 1035
rect -4220 1015 -4200 1035
rect -4130 1015 -4110 1035
rect -4040 1015 -4020 1035
rect -3950 1015 -3930 1035
rect -3860 1015 -3840 1035
rect -3770 1015 -3750 1035
rect -3680 1015 -3660 1035
rect -3590 1015 -3570 1035
rect -3500 1015 -3480 1035
rect -3410 1015 -3390 1035
rect -3320 1015 -3300 1035
rect -3230 1015 -3210 1035
rect -3140 1015 -3120 1035
rect -3050 1015 -3030 1035
rect -2960 1015 -2940 1035
rect -2870 1015 -2850 1035
rect -2780 1015 -2760 1035
rect -2690 1015 -2670 1035
rect -2600 1015 -2580 1035
rect -2510 1015 -2490 1035
rect -2420 1015 -2400 1035
rect -2330 1015 -2310 1035
rect -2240 1015 -2220 1035
rect -2150 1015 -2130 1035
rect -2060 1015 -2040 1035
rect -1970 1015 -1950 1035
rect -1880 1015 -1860 1035
rect -1790 1015 -1770 1035
rect -1700 1015 -1680 1035
rect -1610 1015 -1590 1035
rect -1520 1015 -1500 1035
rect -1430 1015 -1410 1035
rect -1340 1015 -1320 1035
rect -1250 1015 -1230 1035
rect -1160 1015 -1140 1035
rect -1070 1015 -1050 1035
rect -980 1015 -960 1035
rect -890 1015 -870 1035
rect -800 1015 -780 1035
rect -710 1015 -690 1035
rect -620 1015 -600 1035
rect -530 1015 -510 1035
rect -440 1015 -420 1035
rect -350 1015 -330 1035
rect -260 1015 -240 1035
rect -170 1015 -150 1035
rect -80 1015 -60 1035
rect -11510 960 -11490 980
rect -11420 960 -11400 980
rect -11330 960 -11310 980
rect -11240 960 -11220 980
rect -11150 960 -11130 980
rect -11060 960 -11040 980
rect -10970 960 -10950 980
rect -10880 960 -10860 980
rect -10790 960 -10770 980
rect -10700 960 -10680 980
rect -10610 960 -10590 980
rect -10520 960 -10500 980
rect -10430 960 -10410 980
rect -10340 960 -10320 980
rect -10250 960 -10230 980
rect -10160 960 -10140 980
rect -10070 960 -10050 980
rect -9980 960 -9960 980
rect -9890 960 -9870 980
rect -9800 960 -9780 980
rect -9710 960 -9690 980
rect -9620 960 -9600 980
rect -9530 960 -9510 980
rect -9440 960 -9420 980
rect -9350 960 -9330 980
rect -9260 960 -9240 980
rect -9170 960 -9150 980
rect -9080 960 -9060 980
rect -8990 960 -8970 980
rect -8900 960 -8880 980
rect -8810 960 -8790 980
rect -8720 960 -8700 980
rect -8630 960 -8610 980
rect -8540 960 -8520 980
rect -8450 960 -8430 980
rect -8360 960 -8340 980
rect -8270 960 -8250 980
rect -8180 960 -8160 980
rect -8090 960 -8070 980
rect -8000 960 -7980 980
rect -7910 960 -7890 980
rect -7820 960 -7800 980
rect -7730 960 -7710 980
rect -7640 960 -7620 980
rect -7550 960 -7530 980
rect -7460 960 -7440 980
rect -7370 960 -7350 980
rect -7280 960 -7260 980
rect -7190 960 -7170 980
rect -7100 960 -7080 980
rect -7010 960 -6990 980
rect -6920 960 -6900 980
rect -6830 960 -6810 980
rect -6740 960 -6720 980
rect -6650 960 -6630 980
rect -6560 960 -6540 980
rect -6470 960 -6450 980
rect -6380 960 -6360 980
rect -6290 960 -6270 980
rect -6200 960 -6180 980
rect -6110 960 -6090 980
rect -6020 960 -6000 980
rect -5930 960 -5910 980
rect -5840 960 -5820 980
rect -5750 960 -5730 980
rect -5660 960 -5640 980
rect -5570 960 -5550 980
rect -5480 960 -5460 980
rect -5390 960 -5370 980
rect -5300 960 -5280 980
rect -5210 960 -5190 980
rect -5120 960 -5100 980
rect -5030 960 -5010 980
rect -4940 960 -4920 980
rect -4850 960 -4830 980
rect -4760 960 -4740 980
rect -4670 960 -4650 980
rect -4580 960 -4560 980
rect -4490 960 -4470 980
rect -4400 960 -4380 980
rect -4310 960 -4290 980
rect -4220 960 -4200 980
rect -4130 960 -4110 980
rect -4040 960 -4020 980
rect -3950 960 -3930 980
rect -3860 960 -3840 980
rect -3770 960 -3750 980
rect -3680 960 -3660 980
rect -3590 960 -3570 980
rect -3500 960 -3480 980
rect -3410 960 -3390 980
rect -3320 960 -3300 980
rect -3230 960 -3210 980
rect -3140 960 -3120 980
rect -3050 960 -3030 980
rect -2960 960 -2940 980
rect -2870 960 -2850 980
rect -2780 960 -2760 980
rect -2690 960 -2670 980
rect -2600 960 -2580 980
rect -2510 960 -2490 980
rect -2420 960 -2400 980
rect -2330 960 -2310 980
rect -2240 960 -2220 980
rect -2150 960 -2130 980
rect -2060 960 -2040 980
rect -1970 960 -1950 980
rect -1880 960 -1860 980
rect -1790 960 -1770 980
rect -1700 960 -1680 980
rect -1610 960 -1590 980
rect -1520 960 -1500 980
rect -1430 960 -1410 980
rect -1340 960 -1320 980
rect -1250 960 -1230 980
rect -1160 960 -1140 980
rect -1070 960 -1050 980
rect -980 960 -960 980
rect -890 960 -870 980
rect -800 960 -780 980
rect -710 960 -690 980
rect -620 960 -600 980
rect -530 960 -510 980
rect -440 960 -420 980
rect -350 960 -330 980
rect -260 960 -240 980
rect -170 960 -150 980
rect -80 960 -60 980
rect -11510 740 -11490 760
rect -11420 740 -11400 760
rect -11330 740 -11310 760
rect -11240 740 -11220 760
rect -11150 740 -11130 760
rect -11060 740 -11040 760
rect -10970 740 -10950 760
rect -10880 740 -10860 760
rect -10790 740 -10770 760
rect -10700 740 -10680 760
rect -10610 740 -10590 760
rect -10520 740 -10500 760
rect -10430 740 -10410 760
rect -10340 740 -10320 760
rect -10250 740 -10230 760
rect -10160 740 -10140 760
rect -10070 740 -10050 760
rect -9980 740 -9960 760
rect -9890 740 -9870 760
rect -9800 740 -9780 760
rect -9710 740 -9690 760
rect -9620 740 -9600 760
rect -9530 740 -9510 760
rect -9440 740 -9420 760
rect -9350 740 -9330 760
rect -9260 740 -9240 760
rect -9170 740 -9150 760
rect -9080 740 -9060 760
rect -8990 740 -8970 760
rect -8900 740 -8880 760
rect -8810 740 -8790 760
rect -8720 740 -8700 760
rect -8630 740 -8610 760
rect -8540 740 -8520 760
rect -8450 740 -8430 760
rect -8360 740 -8340 760
rect -8270 740 -8250 760
rect -8180 740 -8160 760
rect -8090 740 -8070 760
rect -8000 740 -7980 760
rect -7910 740 -7890 760
rect -7820 740 -7800 760
rect -7730 740 -7710 760
rect -7640 740 -7620 760
rect -7550 740 -7530 760
rect -7460 740 -7440 760
rect -7370 740 -7350 760
rect -7280 740 -7260 760
rect -7190 740 -7170 760
rect -7100 740 -7080 760
rect -7010 740 -6990 760
rect -6920 740 -6900 760
rect -6830 740 -6810 760
rect -6740 740 -6720 760
rect -6650 740 -6630 760
rect -6560 740 -6540 760
rect -6470 740 -6450 760
rect -6380 740 -6360 760
rect -6290 740 -6270 760
rect -6200 740 -6180 760
rect -6110 740 -6090 760
rect -6020 740 -6000 760
rect -5930 740 -5910 760
rect -5840 740 -5820 760
rect -5750 740 -5730 760
rect -5660 740 -5640 760
rect -5570 740 -5550 760
rect -5480 740 -5460 760
rect -5390 740 -5370 760
rect -5300 740 -5280 760
rect -5210 740 -5190 760
rect -5120 740 -5100 760
rect -5030 740 -5010 760
rect -4940 740 -4920 760
rect -4850 740 -4830 760
rect -4760 740 -4740 760
rect -4670 740 -4650 760
rect -4580 740 -4560 760
rect -4490 740 -4470 760
rect -4400 740 -4380 760
rect -4310 740 -4290 760
rect -4220 740 -4200 760
rect -4130 740 -4110 760
rect -4040 740 -4020 760
rect -3950 740 -3930 760
rect -3860 740 -3840 760
rect -3770 740 -3750 760
rect -3680 740 -3660 760
rect -3590 740 -3570 760
rect -3500 740 -3480 760
rect -3410 740 -3390 760
rect -3320 740 -3300 760
rect -3230 740 -3210 760
rect -3140 740 -3120 760
rect -3050 740 -3030 760
rect -2960 740 -2940 760
rect -2870 740 -2850 760
rect -2780 740 -2760 760
rect -2690 740 -2670 760
rect -2600 740 -2580 760
rect -2510 740 -2490 760
rect -2420 740 -2400 760
rect -2330 740 -2310 760
rect -2240 740 -2220 760
rect -2150 740 -2130 760
rect -2060 740 -2040 760
rect -1970 740 -1950 760
rect -1880 740 -1860 760
rect -1790 740 -1770 760
rect -1700 740 -1680 760
rect -1610 740 -1590 760
rect -1520 740 -1500 760
rect -1430 740 -1410 760
rect -1340 740 -1320 760
rect -1250 740 -1230 760
rect -1160 740 -1140 760
rect -1070 740 -1050 760
rect -980 740 -960 760
rect -890 740 -870 760
rect -800 740 -780 760
rect -710 740 -690 760
rect -620 740 -600 760
rect -530 740 -510 760
rect -440 740 -420 760
rect -350 740 -330 760
rect -260 740 -240 760
rect -170 740 -150 760
rect -80 740 -60 760
<< poly >>
rect -11525 1945 -11475 1960
rect -11435 1945 -11385 1960
rect -11345 1945 -11295 1960
rect -11255 1945 -11205 1960
rect -11165 1945 -11115 1960
rect -11075 1945 -11025 1960
rect -10985 1945 -10935 1960
rect -10895 1945 -10845 1960
rect -10805 1945 -10755 1960
rect -10715 1945 -10665 1960
rect -10625 1945 -10575 1960
rect -10535 1945 -10485 1960
rect -10445 1945 -10395 1960
rect -10355 1945 -10305 1960
rect -10265 1945 -10215 1960
rect -10175 1945 -10125 1960
rect -10085 1945 -10035 1960
rect -9995 1945 -9945 1960
rect -9905 1945 -9855 1960
rect -9815 1945 -9765 1960
rect -9725 1945 -9675 1960
rect -9635 1945 -9585 1960
rect -9545 1945 -9495 1960
rect -9455 1945 -9405 1960
rect -9365 1945 -9315 1960
rect -9275 1945 -9225 1960
rect -9185 1945 -9135 1960
rect -9095 1945 -9045 1960
rect -9005 1945 -8955 1960
rect -8915 1945 -8865 1960
rect -8825 1945 -8775 1960
rect -8735 1945 -8685 1960
rect -8645 1945 -8595 1960
rect -8555 1945 -8505 1960
rect -8465 1945 -8415 1960
rect -8375 1945 -8325 1960
rect -8285 1945 -8235 1960
rect -8195 1945 -8145 1960
rect -8105 1945 -8055 1960
rect -8015 1945 -7965 1960
rect -7925 1945 -7875 1960
rect -7835 1945 -7785 1960
rect -7745 1945 -7695 1960
rect -7655 1945 -7605 1960
rect -7565 1945 -7515 1960
rect -7475 1945 -7425 1960
rect -7385 1945 -7335 1960
rect -7295 1945 -7245 1960
rect -7205 1945 -7155 1960
rect -7115 1945 -7065 1960
rect -7025 1945 -6975 1960
rect -6935 1945 -6885 1960
rect -6845 1945 -6795 1960
rect -6755 1945 -6705 1960
rect -6665 1945 -6615 1960
rect -6575 1945 -6525 1960
rect -6485 1945 -6435 1960
rect -6395 1945 -6345 1960
rect -6305 1945 -6255 1960
rect -6215 1945 -6165 1960
rect -6125 1945 -6075 1960
rect -6035 1945 -5985 1960
rect -5945 1945 -5895 1960
rect -5855 1945 -5805 1960
rect -5765 1945 -5715 1960
rect -5675 1945 -5625 1960
rect -5585 1945 -5535 1960
rect -5495 1945 -5445 1960
rect -5405 1945 -5355 1960
rect -5315 1945 -5265 1960
rect -5225 1945 -5175 1960
rect -5135 1945 -5085 1960
rect -5045 1945 -4995 1960
rect -4955 1945 -4905 1960
rect -4865 1945 -4815 1960
rect -4775 1945 -4725 1960
rect -4685 1945 -4635 1960
rect -4595 1945 -4545 1960
rect -4505 1945 -4455 1960
rect -4415 1945 -4365 1960
rect -4325 1945 -4275 1960
rect -4235 1945 -4185 1960
rect -4145 1945 -4095 1960
rect -4055 1945 -4005 1960
rect -3965 1945 -3915 1960
rect -3875 1945 -3825 1960
rect -3785 1945 -3735 1960
rect -3695 1945 -3645 1960
rect -3605 1945 -3555 1960
rect -3515 1945 -3465 1960
rect -3425 1945 -3375 1960
rect -3335 1945 -3285 1960
rect -3245 1945 -3195 1960
rect -3155 1945 -3105 1960
rect -3065 1945 -3015 1960
rect -2975 1945 -2925 1960
rect -2885 1945 -2835 1960
rect -2795 1945 -2745 1960
rect -2705 1945 -2655 1960
rect -2615 1945 -2565 1960
rect -2525 1945 -2475 1960
rect -2435 1945 -2385 1960
rect -2345 1945 -2295 1960
rect -2255 1945 -2205 1960
rect -2165 1945 -2115 1960
rect -2075 1945 -2025 1960
rect -1985 1945 -1935 1960
rect -1895 1945 -1845 1960
rect -1805 1945 -1755 1960
rect -1715 1945 -1665 1960
rect -1625 1945 -1575 1960
rect -1535 1945 -1485 1960
rect -1445 1945 -1395 1960
rect -1355 1945 -1305 1960
rect -1265 1945 -1215 1960
rect -1175 1945 -1125 1960
rect -1085 1945 -1035 1960
rect -995 1945 -945 1960
rect -905 1945 -855 1960
rect -815 1945 -765 1960
rect -725 1945 -675 1960
rect -635 1945 -585 1960
rect -545 1945 -495 1960
rect -455 1945 -405 1960
rect -365 1945 -315 1960
rect -275 1945 -225 1960
rect -185 1945 -135 1960
rect -95 1945 -45 1960
rect -11525 1825 -11475 1845
rect -11435 1825 -11385 1845
rect -11525 1820 -11385 1825
rect -11525 1800 -11510 1820
rect -11490 1800 -11420 1820
rect -11400 1800 -11385 1820
rect -11525 1795 -11385 1800
rect -11345 1825 -11295 1845
rect -11255 1825 -11205 1845
rect -11345 1820 -11205 1825
rect -11345 1800 -11330 1820
rect -11310 1800 -11240 1820
rect -11220 1800 -11205 1820
rect -11345 1795 -11205 1800
rect -11165 1825 -11115 1845
rect -11075 1825 -11025 1845
rect -11165 1820 -11025 1825
rect -11165 1800 -11150 1820
rect -11130 1800 -11060 1820
rect -11040 1800 -11025 1820
rect -11165 1795 -11025 1800
rect -10985 1825 -10935 1845
rect -10895 1825 -10845 1845
rect -10985 1820 -10845 1825
rect -10985 1800 -10970 1820
rect -10950 1800 -10880 1820
rect -10860 1800 -10845 1820
rect -10985 1795 -10845 1800
rect -10805 1825 -10755 1845
rect -10715 1825 -10665 1845
rect -10805 1820 -10665 1825
rect -10805 1800 -10790 1820
rect -10770 1800 -10700 1820
rect -10680 1800 -10665 1820
rect -10805 1795 -10665 1800
rect -10625 1825 -10575 1845
rect -10535 1825 -10485 1845
rect -10625 1820 -10485 1825
rect -10625 1800 -10610 1820
rect -10590 1800 -10520 1820
rect -10500 1800 -10485 1820
rect -10625 1795 -10485 1800
rect -10445 1825 -10395 1845
rect -10355 1825 -10305 1845
rect -10445 1820 -10305 1825
rect -10445 1800 -10430 1820
rect -10410 1800 -10340 1820
rect -10320 1800 -10305 1820
rect -10445 1795 -10305 1800
rect -10265 1825 -10215 1845
rect -10175 1825 -10125 1845
rect -10265 1820 -10125 1825
rect -10265 1800 -10250 1820
rect -10230 1800 -10160 1820
rect -10140 1800 -10125 1820
rect -10265 1795 -10125 1800
rect -10085 1825 -10035 1845
rect -9995 1825 -9945 1845
rect -10085 1820 -9945 1825
rect -10085 1800 -10070 1820
rect -10050 1800 -9980 1820
rect -9960 1800 -9945 1820
rect -10085 1795 -9945 1800
rect -9905 1825 -9855 1845
rect -9815 1825 -9765 1845
rect -9905 1820 -9765 1825
rect -9905 1800 -9890 1820
rect -9870 1800 -9800 1820
rect -9780 1800 -9765 1820
rect -9905 1795 -9765 1800
rect -9725 1825 -9675 1845
rect -9635 1825 -9585 1845
rect -9725 1820 -9585 1825
rect -9725 1800 -9710 1820
rect -9690 1800 -9620 1820
rect -9600 1800 -9585 1820
rect -9725 1795 -9585 1800
rect -9545 1825 -9495 1845
rect -9455 1825 -9405 1845
rect -9545 1820 -9405 1825
rect -9545 1800 -9530 1820
rect -9510 1800 -9440 1820
rect -9420 1800 -9405 1820
rect -9545 1795 -9405 1800
rect -9365 1825 -9315 1845
rect -9275 1825 -9225 1845
rect -9365 1820 -9225 1825
rect -9365 1800 -9350 1820
rect -9330 1800 -9260 1820
rect -9240 1800 -9225 1820
rect -9365 1795 -9225 1800
rect -9185 1825 -9135 1845
rect -9095 1825 -9045 1845
rect -9185 1820 -9045 1825
rect -9185 1800 -9170 1820
rect -9150 1800 -9080 1820
rect -9060 1800 -9045 1820
rect -9185 1795 -9045 1800
rect -9005 1825 -8955 1845
rect -8915 1825 -8865 1845
rect -9005 1820 -8865 1825
rect -9005 1800 -8990 1820
rect -8970 1800 -8900 1820
rect -8880 1800 -8865 1820
rect -9005 1795 -8865 1800
rect -8825 1825 -8775 1845
rect -8735 1825 -8685 1845
rect -8825 1820 -8685 1825
rect -8825 1800 -8810 1820
rect -8790 1800 -8720 1820
rect -8700 1800 -8685 1820
rect -8825 1795 -8685 1800
rect -8645 1825 -8595 1845
rect -8555 1825 -8505 1845
rect -8645 1820 -8505 1825
rect -8645 1800 -8630 1820
rect -8610 1800 -8540 1820
rect -8520 1800 -8505 1820
rect -8645 1795 -8505 1800
rect -8465 1825 -8415 1845
rect -8375 1825 -8325 1845
rect -8465 1820 -8325 1825
rect -8465 1800 -8450 1820
rect -8430 1800 -8360 1820
rect -8340 1800 -8325 1820
rect -8465 1795 -8325 1800
rect -8285 1825 -8235 1845
rect -8195 1825 -8145 1845
rect -8285 1820 -8145 1825
rect -8285 1800 -8270 1820
rect -8250 1800 -8180 1820
rect -8160 1800 -8145 1820
rect -8285 1795 -8145 1800
rect -8105 1825 -8055 1845
rect -8015 1825 -7965 1845
rect -8105 1820 -7965 1825
rect -8105 1800 -8090 1820
rect -8070 1800 -8000 1820
rect -7980 1800 -7965 1820
rect -8105 1795 -7965 1800
rect -7925 1825 -7875 1845
rect -7835 1825 -7785 1845
rect -7925 1820 -7785 1825
rect -7925 1800 -7910 1820
rect -7890 1800 -7820 1820
rect -7800 1800 -7785 1820
rect -7925 1795 -7785 1800
rect -7745 1825 -7695 1845
rect -7655 1825 -7605 1845
rect -7745 1820 -7605 1825
rect -7745 1800 -7730 1820
rect -7710 1800 -7640 1820
rect -7620 1800 -7605 1820
rect -7745 1795 -7605 1800
rect -7565 1825 -7515 1845
rect -7475 1825 -7425 1845
rect -7565 1820 -7425 1825
rect -7565 1800 -7550 1820
rect -7530 1800 -7460 1820
rect -7440 1800 -7425 1820
rect -7565 1795 -7425 1800
rect -7385 1825 -7335 1845
rect -7295 1825 -7245 1845
rect -7385 1820 -7245 1825
rect -7385 1800 -7370 1820
rect -7350 1800 -7280 1820
rect -7260 1800 -7245 1820
rect -7385 1795 -7245 1800
rect -7205 1825 -7155 1845
rect -7115 1825 -7065 1845
rect -7205 1820 -7065 1825
rect -7205 1800 -7190 1820
rect -7170 1800 -7100 1820
rect -7080 1800 -7065 1820
rect -7205 1795 -7065 1800
rect -7025 1825 -6975 1845
rect -6935 1825 -6885 1845
rect -7025 1820 -6885 1825
rect -7025 1800 -7010 1820
rect -6990 1800 -6920 1820
rect -6900 1800 -6885 1820
rect -7025 1795 -6885 1800
rect -6845 1825 -6795 1845
rect -6755 1825 -6705 1845
rect -6845 1820 -6705 1825
rect -6845 1800 -6830 1820
rect -6810 1800 -6740 1820
rect -6720 1800 -6705 1820
rect -6845 1795 -6705 1800
rect -6665 1825 -6615 1845
rect -6575 1825 -6525 1845
rect -6665 1820 -6525 1825
rect -6665 1800 -6650 1820
rect -6630 1800 -6560 1820
rect -6540 1800 -6525 1820
rect -6665 1795 -6525 1800
rect -6485 1825 -6435 1845
rect -6395 1825 -6345 1845
rect -6485 1820 -6345 1825
rect -6485 1800 -6470 1820
rect -6450 1800 -6380 1820
rect -6360 1800 -6345 1820
rect -6485 1795 -6345 1800
rect -6305 1825 -6255 1845
rect -6215 1825 -6165 1845
rect -6305 1820 -6165 1825
rect -6305 1800 -6290 1820
rect -6270 1800 -6200 1820
rect -6180 1800 -6165 1820
rect -6305 1795 -6165 1800
rect -6125 1825 -6075 1845
rect -6035 1825 -5985 1845
rect -6125 1820 -5985 1825
rect -6125 1800 -6110 1820
rect -6090 1800 -6020 1820
rect -6000 1800 -5985 1820
rect -6125 1795 -5985 1800
rect -5945 1825 -5895 1845
rect -5855 1825 -5805 1845
rect -5945 1820 -5805 1825
rect -5945 1800 -5930 1820
rect -5910 1800 -5840 1820
rect -5820 1800 -5805 1820
rect -5945 1795 -5805 1800
rect -5765 1825 -5715 1845
rect -5675 1825 -5625 1845
rect -5765 1820 -5625 1825
rect -5765 1800 -5750 1820
rect -5730 1800 -5660 1820
rect -5640 1800 -5625 1820
rect -5765 1795 -5625 1800
rect -5585 1825 -5535 1845
rect -5495 1825 -5445 1845
rect -5585 1820 -5445 1825
rect -5585 1800 -5570 1820
rect -5550 1800 -5480 1820
rect -5460 1800 -5445 1820
rect -5585 1795 -5445 1800
rect -5405 1825 -5355 1845
rect -5315 1825 -5265 1845
rect -5405 1820 -5265 1825
rect -5405 1800 -5390 1820
rect -5370 1800 -5300 1820
rect -5280 1800 -5265 1820
rect -5405 1795 -5265 1800
rect -5225 1825 -5175 1845
rect -5135 1825 -5085 1845
rect -5225 1820 -5085 1825
rect -5225 1800 -5210 1820
rect -5190 1800 -5120 1820
rect -5100 1800 -5085 1820
rect -5225 1795 -5085 1800
rect -5045 1825 -4995 1845
rect -4955 1825 -4905 1845
rect -5045 1820 -4905 1825
rect -5045 1800 -5030 1820
rect -5010 1800 -4940 1820
rect -4920 1800 -4905 1820
rect -5045 1795 -4905 1800
rect -4865 1825 -4815 1845
rect -4775 1825 -4725 1845
rect -4865 1820 -4725 1825
rect -4865 1800 -4850 1820
rect -4830 1800 -4760 1820
rect -4740 1800 -4725 1820
rect -4865 1795 -4725 1800
rect -4685 1825 -4635 1845
rect -4595 1825 -4545 1845
rect -4685 1820 -4545 1825
rect -4685 1800 -4670 1820
rect -4650 1800 -4580 1820
rect -4560 1800 -4545 1820
rect -4685 1795 -4545 1800
rect -4505 1825 -4455 1845
rect -4415 1825 -4365 1845
rect -4505 1820 -4365 1825
rect -4505 1800 -4490 1820
rect -4470 1800 -4400 1820
rect -4380 1800 -4365 1820
rect -4505 1795 -4365 1800
rect -4325 1825 -4275 1845
rect -4235 1825 -4185 1845
rect -4325 1820 -4185 1825
rect -4325 1800 -4310 1820
rect -4290 1800 -4220 1820
rect -4200 1800 -4185 1820
rect -4325 1795 -4185 1800
rect -4145 1825 -4095 1845
rect -4055 1825 -4005 1845
rect -4145 1820 -4005 1825
rect -4145 1800 -4130 1820
rect -4110 1800 -4040 1820
rect -4020 1800 -4005 1820
rect -4145 1795 -4005 1800
rect -3965 1825 -3915 1845
rect -3875 1825 -3825 1845
rect -3965 1820 -3825 1825
rect -3965 1800 -3950 1820
rect -3930 1800 -3860 1820
rect -3840 1800 -3825 1820
rect -3965 1795 -3825 1800
rect -3785 1825 -3735 1845
rect -3695 1825 -3645 1845
rect -3785 1820 -3645 1825
rect -3785 1800 -3770 1820
rect -3750 1800 -3680 1820
rect -3660 1800 -3645 1820
rect -3785 1795 -3645 1800
rect -3605 1825 -3555 1845
rect -3515 1825 -3465 1845
rect -3605 1820 -3465 1825
rect -3605 1800 -3590 1820
rect -3570 1800 -3500 1820
rect -3480 1800 -3465 1820
rect -3605 1795 -3465 1800
rect -3425 1825 -3375 1845
rect -3335 1825 -3285 1845
rect -3425 1820 -3285 1825
rect -3425 1800 -3410 1820
rect -3390 1800 -3320 1820
rect -3300 1800 -3285 1820
rect -3425 1795 -3285 1800
rect -3245 1825 -3195 1845
rect -3155 1825 -3105 1845
rect -3245 1820 -3105 1825
rect -3245 1800 -3230 1820
rect -3210 1800 -3140 1820
rect -3120 1800 -3105 1820
rect -3245 1795 -3105 1800
rect -3065 1825 -3015 1845
rect -2975 1825 -2925 1845
rect -3065 1820 -2925 1825
rect -3065 1800 -3050 1820
rect -3030 1800 -2960 1820
rect -2940 1800 -2925 1820
rect -3065 1795 -2925 1800
rect -2885 1825 -2835 1845
rect -2795 1825 -2745 1845
rect -2885 1820 -2745 1825
rect -2885 1800 -2870 1820
rect -2850 1800 -2780 1820
rect -2760 1800 -2745 1820
rect -2885 1795 -2745 1800
rect -2705 1825 -2655 1845
rect -2615 1825 -2565 1845
rect -2705 1820 -2565 1825
rect -2705 1800 -2690 1820
rect -2670 1800 -2600 1820
rect -2580 1800 -2565 1820
rect -2705 1795 -2565 1800
rect -2525 1825 -2475 1845
rect -2435 1825 -2385 1845
rect -2525 1820 -2385 1825
rect -2525 1800 -2510 1820
rect -2490 1800 -2420 1820
rect -2400 1800 -2385 1820
rect -2525 1795 -2385 1800
rect -2345 1825 -2295 1845
rect -2255 1825 -2205 1845
rect -2345 1820 -2205 1825
rect -2345 1800 -2330 1820
rect -2310 1800 -2240 1820
rect -2220 1800 -2205 1820
rect -2345 1795 -2205 1800
rect -2165 1825 -2115 1845
rect -2075 1825 -2025 1845
rect -2165 1820 -2025 1825
rect -2165 1800 -2150 1820
rect -2130 1800 -2060 1820
rect -2040 1800 -2025 1820
rect -2165 1795 -2025 1800
rect -1985 1825 -1935 1845
rect -1895 1825 -1845 1845
rect -1985 1820 -1845 1825
rect -1985 1800 -1970 1820
rect -1950 1800 -1880 1820
rect -1860 1800 -1845 1820
rect -1985 1795 -1845 1800
rect -1805 1825 -1755 1845
rect -1715 1825 -1665 1845
rect -1805 1820 -1665 1825
rect -1805 1800 -1790 1820
rect -1770 1800 -1700 1820
rect -1680 1800 -1665 1820
rect -1805 1795 -1665 1800
rect -1625 1825 -1575 1845
rect -1535 1825 -1485 1845
rect -1625 1820 -1485 1825
rect -1625 1800 -1610 1820
rect -1590 1800 -1520 1820
rect -1500 1800 -1485 1820
rect -1625 1795 -1485 1800
rect -1445 1825 -1395 1845
rect -1355 1825 -1305 1845
rect -1445 1820 -1305 1825
rect -1445 1800 -1430 1820
rect -1410 1800 -1340 1820
rect -1320 1800 -1305 1820
rect -1445 1795 -1305 1800
rect -1265 1825 -1215 1845
rect -1175 1825 -1125 1845
rect -1265 1820 -1125 1825
rect -1265 1800 -1250 1820
rect -1230 1800 -1160 1820
rect -1140 1800 -1125 1820
rect -1265 1795 -1125 1800
rect -1085 1825 -1035 1845
rect -995 1825 -945 1845
rect -1085 1820 -945 1825
rect -1085 1800 -1070 1820
rect -1050 1800 -980 1820
rect -960 1800 -945 1820
rect -1085 1795 -945 1800
rect -905 1825 -855 1845
rect -815 1825 -765 1845
rect -905 1820 -765 1825
rect -905 1800 -890 1820
rect -870 1800 -800 1820
rect -780 1800 -765 1820
rect -905 1795 -765 1800
rect -725 1825 -675 1845
rect -635 1825 -585 1845
rect -725 1820 -585 1825
rect -725 1800 -710 1820
rect -690 1800 -620 1820
rect -600 1800 -585 1820
rect -725 1795 -585 1800
rect -545 1825 -495 1845
rect -455 1825 -405 1845
rect -545 1820 -405 1825
rect -545 1800 -530 1820
rect -510 1800 -440 1820
rect -420 1800 -405 1820
rect -545 1795 -405 1800
rect -365 1825 -315 1845
rect -275 1825 -225 1845
rect -365 1820 -225 1825
rect -365 1800 -350 1820
rect -330 1800 -260 1820
rect -240 1800 -225 1820
rect -365 1795 -225 1800
rect -185 1825 -135 1845
rect -95 1825 -45 1845
rect -185 1820 -45 1825
rect -185 1800 -170 1820
rect -150 1800 -80 1820
rect -60 1800 -45 1820
rect -185 1795 -45 1800
rect -11525 1210 -11385 1215
rect -11525 1190 -11510 1210
rect -11490 1190 -11420 1210
rect -11400 1190 -11385 1210
rect -11525 1185 -11385 1190
rect -11525 1165 -11475 1185
rect -11435 1165 -11385 1185
rect -11345 1210 -11205 1215
rect -11345 1190 -11330 1210
rect -11310 1190 -11240 1210
rect -11220 1190 -11205 1210
rect -11345 1185 -11205 1190
rect -11345 1165 -11295 1185
rect -11255 1165 -11205 1185
rect -11165 1210 -11025 1215
rect -11165 1190 -11150 1210
rect -11130 1190 -11060 1210
rect -11040 1190 -11025 1210
rect -11165 1185 -11025 1190
rect -11165 1165 -11115 1185
rect -11075 1165 -11025 1185
rect -10985 1210 -10845 1215
rect -10985 1190 -10970 1210
rect -10950 1190 -10880 1210
rect -10860 1190 -10845 1210
rect -10985 1185 -10845 1190
rect -10985 1165 -10935 1185
rect -10895 1165 -10845 1185
rect -10805 1210 -10665 1215
rect -10805 1190 -10790 1210
rect -10770 1190 -10700 1210
rect -10680 1190 -10665 1210
rect -10805 1185 -10665 1190
rect -10805 1165 -10755 1185
rect -10715 1165 -10665 1185
rect -10625 1210 -10485 1215
rect -10625 1190 -10610 1210
rect -10590 1190 -10520 1210
rect -10500 1190 -10485 1210
rect -10625 1185 -10485 1190
rect -10625 1165 -10575 1185
rect -10535 1165 -10485 1185
rect -10445 1210 -10305 1215
rect -10445 1190 -10430 1210
rect -10410 1190 -10340 1210
rect -10320 1190 -10305 1210
rect -10445 1185 -10305 1190
rect -10445 1165 -10395 1185
rect -10355 1165 -10305 1185
rect -10265 1210 -10125 1215
rect -10265 1190 -10250 1210
rect -10230 1190 -10160 1210
rect -10140 1190 -10125 1210
rect -10265 1185 -10125 1190
rect -10265 1165 -10215 1185
rect -10175 1165 -10125 1185
rect -10085 1210 -9945 1215
rect -10085 1190 -10070 1210
rect -10050 1190 -9980 1210
rect -9960 1190 -9945 1210
rect -10085 1185 -9945 1190
rect -10085 1165 -10035 1185
rect -9995 1165 -9945 1185
rect -9905 1210 -9765 1215
rect -9905 1190 -9890 1210
rect -9870 1190 -9800 1210
rect -9780 1190 -9765 1210
rect -9905 1185 -9765 1190
rect -9905 1165 -9855 1185
rect -9815 1165 -9765 1185
rect -9725 1210 -9585 1215
rect -9725 1190 -9710 1210
rect -9690 1190 -9620 1210
rect -9600 1190 -9585 1210
rect -9725 1185 -9585 1190
rect -9725 1165 -9675 1185
rect -9635 1165 -9585 1185
rect -9545 1210 -9405 1215
rect -9545 1190 -9530 1210
rect -9510 1190 -9440 1210
rect -9420 1190 -9405 1210
rect -9545 1185 -9405 1190
rect -9545 1165 -9495 1185
rect -9455 1165 -9405 1185
rect -9365 1210 -9225 1215
rect -9365 1190 -9350 1210
rect -9330 1190 -9260 1210
rect -9240 1190 -9225 1210
rect -9365 1185 -9225 1190
rect -9365 1165 -9315 1185
rect -9275 1165 -9225 1185
rect -9185 1210 -9045 1215
rect -9185 1190 -9170 1210
rect -9150 1190 -9080 1210
rect -9060 1190 -9045 1210
rect -9185 1185 -9045 1190
rect -9185 1165 -9135 1185
rect -9095 1165 -9045 1185
rect -9005 1210 -8865 1215
rect -9005 1190 -8990 1210
rect -8970 1190 -8900 1210
rect -8880 1190 -8865 1210
rect -9005 1185 -8865 1190
rect -9005 1165 -8955 1185
rect -8915 1165 -8865 1185
rect -8825 1210 -8685 1215
rect -8825 1190 -8810 1210
rect -8790 1190 -8720 1210
rect -8700 1190 -8685 1210
rect -8825 1185 -8685 1190
rect -8825 1165 -8775 1185
rect -8735 1165 -8685 1185
rect -8645 1210 -8505 1215
rect -8645 1190 -8630 1210
rect -8610 1190 -8540 1210
rect -8520 1190 -8505 1210
rect -8645 1185 -8505 1190
rect -8645 1165 -8595 1185
rect -8555 1165 -8505 1185
rect -8465 1210 -8325 1215
rect -8465 1190 -8450 1210
rect -8430 1190 -8360 1210
rect -8340 1190 -8325 1210
rect -8465 1185 -8325 1190
rect -8465 1165 -8415 1185
rect -8375 1165 -8325 1185
rect -8285 1210 -8145 1215
rect -8285 1190 -8270 1210
rect -8250 1190 -8180 1210
rect -8160 1190 -8145 1210
rect -8285 1185 -8145 1190
rect -8285 1165 -8235 1185
rect -8195 1165 -8145 1185
rect -8105 1210 -7965 1215
rect -8105 1190 -8090 1210
rect -8070 1190 -8000 1210
rect -7980 1190 -7965 1210
rect -8105 1185 -7965 1190
rect -8105 1165 -8055 1185
rect -8015 1165 -7965 1185
rect -7925 1210 -7785 1215
rect -7925 1190 -7910 1210
rect -7890 1190 -7820 1210
rect -7800 1190 -7785 1210
rect -7925 1185 -7785 1190
rect -7925 1165 -7875 1185
rect -7835 1165 -7785 1185
rect -7745 1210 -7605 1215
rect -7745 1190 -7730 1210
rect -7710 1190 -7640 1210
rect -7620 1190 -7605 1210
rect -7745 1185 -7605 1190
rect -7745 1165 -7695 1185
rect -7655 1165 -7605 1185
rect -7565 1210 -7425 1215
rect -7565 1190 -7550 1210
rect -7530 1190 -7460 1210
rect -7440 1190 -7425 1210
rect -7565 1185 -7425 1190
rect -7565 1165 -7515 1185
rect -7475 1165 -7425 1185
rect -7385 1210 -7245 1215
rect -7385 1190 -7370 1210
rect -7350 1190 -7280 1210
rect -7260 1190 -7245 1210
rect -7385 1185 -7245 1190
rect -7385 1165 -7335 1185
rect -7295 1165 -7245 1185
rect -7205 1210 -7065 1215
rect -7205 1190 -7190 1210
rect -7170 1190 -7100 1210
rect -7080 1190 -7065 1210
rect -7205 1185 -7065 1190
rect -7205 1165 -7155 1185
rect -7115 1165 -7065 1185
rect -7025 1210 -6885 1215
rect -7025 1190 -7010 1210
rect -6990 1190 -6920 1210
rect -6900 1190 -6885 1210
rect -7025 1185 -6885 1190
rect -7025 1165 -6975 1185
rect -6935 1165 -6885 1185
rect -6845 1210 -6705 1215
rect -6845 1190 -6830 1210
rect -6810 1190 -6740 1210
rect -6720 1190 -6705 1210
rect -6845 1185 -6705 1190
rect -6845 1165 -6795 1185
rect -6755 1165 -6705 1185
rect -6665 1210 -6525 1215
rect -6665 1190 -6650 1210
rect -6630 1190 -6560 1210
rect -6540 1190 -6525 1210
rect -6665 1185 -6525 1190
rect -6665 1165 -6615 1185
rect -6575 1165 -6525 1185
rect -6485 1210 -6345 1215
rect -6485 1190 -6470 1210
rect -6450 1190 -6380 1210
rect -6360 1190 -6345 1210
rect -6485 1185 -6345 1190
rect -6485 1165 -6435 1185
rect -6395 1165 -6345 1185
rect -6305 1210 -6165 1215
rect -6305 1190 -6290 1210
rect -6270 1190 -6200 1210
rect -6180 1190 -6165 1210
rect -6305 1185 -6165 1190
rect -6305 1165 -6255 1185
rect -6215 1165 -6165 1185
rect -6125 1210 -5985 1215
rect -6125 1190 -6110 1210
rect -6090 1190 -6020 1210
rect -6000 1190 -5985 1210
rect -6125 1185 -5985 1190
rect -6125 1165 -6075 1185
rect -6035 1165 -5985 1185
rect -5945 1210 -5805 1215
rect -5945 1190 -5930 1210
rect -5910 1190 -5840 1210
rect -5820 1190 -5805 1210
rect -5945 1185 -5805 1190
rect -5945 1165 -5895 1185
rect -5855 1165 -5805 1185
rect -5765 1210 -5625 1215
rect -5765 1190 -5750 1210
rect -5730 1190 -5660 1210
rect -5640 1190 -5625 1210
rect -5765 1185 -5625 1190
rect -5765 1165 -5715 1185
rect -5675 1165 -5625 1185
rect -5585 1210 -5445 1215
rect -5585 1190 -5570 1210
rect -5550 1190 -5480 1210
rect -5460 1190 -5445 1210
rect -5585 1185 -5445 1190
rect -5585 1165 -5535 1185
rect -5495 1165 -5445 1185
rect -5405 1210 -5265 1215
rect -5405 1190 -5390 1210
rect -5370 1190 -5300 1210
rect -5280 1190 -5265 1210
rect -5405 1185 -5265 1190
rect -5405 1165 -5355 1185
rect -5315 1165 -5265 1185
rect -5225 1210 -5085 1215
rect -5225 1190 -5210 1210
rect -5190 1190 -5120 1210
rect -5100 1190 -5085 1210
rect -5225 1185 -5085 1190
rect -5225 1165 -5175 1185
rect -5135 1165 -5085 1185
rect -5045 1210 -4905 1215
rect -5045 1190 -5030 1210
rect -5010 1190 -4940 1210
rect -4920 1190 -4905 1210
rect -5045 1185 -4905 1190
rect -5045 1165 -4995 1185
rect -4955 1165 -4905 1185
rect -4865 1210 -4725 1215
rect -4865 1190 -4850 1210
rect -4830 1190 -4760 1210
rect -4740 1190 -4725 1210
rect -4865 1185 -4725 1190
rect -4865 1165 -4815 1185
rect -4775 1165 -4725 1185
rect -4685 1210 -4545 1215
rect -4685 1190 -4670 1210
rect -4650 1190 -4580 1210
rect -4560 1190 -4545 1210
rect -4685 1185 -4545 1190
rect -4685 1165 -4635 1185
rect -4595 1165 -4545 1185
rect -4505 1210 -4365 1215
rect -4505 1190 -4490 1210
rect -4470 1190 -4400 1210
rect -4380 1190 -4365 1210
rect -4505 1185 -4365 1190
rect -4505 1165 -4455 1185
rect -4415 1165 -4365 1185
rect -4325 1210 -4185 1215
rect -4325 1190 -4310 1210
rect -4290 1190 -4220 1210
rect -4200 1190 -4185 1210
rect -4325 1185 -4185 1190
rect -4325 1165 -4275 1185
rect -4235 1165 -4185 1185
rect -4145 1210 -4005 1215
rect -4145 1190 -4130 1210
rect -4110 1190 -4040 1210
rect -4020 1190 -4005 1210
rect -4145 1185 -4005 1190
rect -4145 1165 -4095 1185
rect -4055 1165 -4005 1185
rect -3965 1210 -3825 1215
rect -3965 1190 -3950 1210
rect -3930 1190 -3860 1210
rect -3840 1190 -3825 1210
rect -3965 1185 -3825 1190
rect -3965 1165 -3915 1185
rect -3875 1165 -3825 1185
rect -3785 1210 -3645 1215
rect -3785 1190 -3770 1210
rect -3750 1190 -3680 1210
rect -3660 1190 -3645 1210
rect -3785 1185 -3645 1190
rect -3785 1165 -3735 1185
rect -3695 1165 -3645 1185
rect -3605 1210 -3465 1215
rect -3605 1190 -3590 1210
rect -3570 1190 -3500 1210
rect -3480 1190 -3465 1210
rect -3605 1185 -3465 1190
rect -3605 1165 -3555 1185
rect -3515 1165 -3465 1185
rect -3425 1210 -3285 1215
rect -3425 1190 -3410 1210
rect -3390 1190 -3320 1210
rect -3300 1190 -3285 1210
rect -3425 1185 -3285 1190
rect -3425 1165 -3375 1185
rect -3335 1165 -3285 1185
rect -3245 1210 -3105 1215
rect -3245 1190 -3230 1210
rect -3210 1190 -3140 1210
rect -3120 1190 -3105 1210
rect -3245 1185 -3105 1190
rect -3245 1165 -3195 1185
rect -3155 1165 -3105 1185
rect -3065 1210 -2925 1215
rect -3065 1190 -3050 1210
rect -3030 1190 -2960 1210
rect -2940 1190 -2925 1210
rect -3065 1185 -2925 1190
rect -3065 1165 -3015 1185
rect -2975 1165 -2925 1185
rect -2885 1210 -2745 1215
rect -2885 1190 -2870 1210
rect -2850 1190 -2780 1210
rect -2760 1190 -2745 1210
rect -2885 1185 -2745 1190
rect -2885 1165 -2835 1185
rect -2795 1165 -2745 1185
rect -2705 1210 -2565 1215
rect -2705 1190 -2690 1210
rect -2670 1190 -2600 1210
rect -2580 1190 -2565 1210
rect -2705 1185 -2565 1190
rect -2705 1165 -2655 1185
rect -2615 1165 -2565 1185
rect -2525 1210 -2385 1215
rect -2525 1190 -2510 1210
rect -2490 1190 -2420 1210
rect -2400 1190 -2385 1210
rect -2525 1185 -2385 1190
rect -2525 1165 -2475 1185
rect -2435 1165 -2385 1185
rect -2345 1210 -2205 1215
rect -2345 1190 -2330 1210
rect -2310 1190 -2240 1210
rect -2220 1190 -2205 1210
rect -2345 1185 -2205 1190
rect -2345 1165 -2295 1185
rect -2255 1165 -2205 1185
rect -2165 1210 -2025 1215
rect -2165 1190 -2150 1210
rect -2130 1190 -2060 1210
rect -2040 1190 -2025 1210
rect -2165 1185 -2025 1190
rect -2165 1165 -2115 1185
rect -2075 1165 -2025 1185
rect -1985 1210 -1845 1215
rect -1985 1190 -1970 1210
rect -1950 1190 -1880 1210
rect -1860 1190 -1845 1210
rect -1985 1185 -1845 1190
rect -1985 1165 -1935 1185
rect -1895 1165 -1845 1185
rect -1805 1210 -1665 1215
rect -1805 1190 -1790 1210
rect -1770 1190 -1700 1210
rect -1680 1190 -1665 1210
rect -1805 1185 -1665 1190
rect -1805 1165 -1755 1185
rect -1715 1165 -1665 1185
rect -1625 1210 -1485 1215
rect -1625 1190 -1610 1210
rect -1590 1190 -1520 1210
rect -1500 1190 -1485 1210
rect -1625 1185 -1485 1190
rect -1625 1165 -1575 1185
rect -1535 1165 -1485 1185
rect -1445 1210 -1305 1215
rect -1445 1190 -1430 1210
rect -1410 1190 -1340 1210
rect -1320 1190 -1305 1210
rect -1445 1185 -1305 1190
rect -1445 1165 -1395 1185
rect -1355 1165 -1305 1185
rect -1265 1210 -1125 1215
rect -1265 1190 -1250 1210
rect -1230 1190 -1160 1210
rect -1140 1190 -1125 1210
rect -1265 1185 -1125 1190
rect -1265 1165 -1215 1185
rect -1175 1165 -1125 1185
rect -1085 1210 -945 1215
rect -1085 1190 -1070 1210
rect -1050 1190 -980 1210
rect -960 1190 -945 1210
rect -1085 1185 -945 1190
rect -1085 1165 -1035 1185
rect -995 1165 -945 1185
rect -905 1210 -765 1215
rect -905 1190 -890 1210
rect -870 1190 -800 1210
rect -780 1190 -765 1210
rect -905 1185 -765 1190
rect -905 1165 -855 1185
rect -815 1165 -765 1185
rect -725 1210 -585 1215
rect -725 1190 -710 1210
rect -690 1190 -620 1210
rect -600 1190 -585 1210
rect -725 1185 -585 1190
rect -725 1165 -675 1185
rect -635 1165 -585 1185
rect -545 1210 -405 1215
rect -545 1190 -530 1210
rect -510 1190 -440 1210
rect -420 1190 -405 1210
rect -545 1185 -405 1190
rect -545 1165 -495 1185
rect -455 1165 -405 1185
rect -365 1210 -225 1215
rect -365 1190 -350 1210
rect -330 1190 -260 1210
rect -240 1190 -225 1210
rect -365 1185 -225 1190
rect -365 1165 -315 1185
rect -275 1165 -225 1185
rect -185 1210 -45 1215
rect -185 1190 -170 1210
rect -150 1190 -80 1210
rect -60 1190 -45 1210
rect -185 1185 -45 1190
rect -185 1165 -135 1185
rect -95 1165 -45 1185
rect -11525 1050 -11475 1065
rect -11435 1050 -11385 1065
rect -11345 1050 -11295 1065
rect -11255 1050 -11205 1065
rect -11165 1050 -11115 1065
rect -11075 1050 -11025 1065
rect -10985 1050 -10935 1065
rect -10895 1050 -10845 1065
rect -10805 1050 -10755 1065
rect -10715 1050 -10665 1065
rect -10625 1050 -10575 1065
rect -10535 1050 -10485 1065
rect -10445 1050 -10395 1065
rect -10355 1050 -10305 1065
rect -10265 1050 -10215 1065
rect -10175 1050 -10125 1065
rect -10085 1050 -10035 1065
rect -9995 1050 -9945 1065
rect -9905 1050 -9855 1065
rect -9815 1050 -9765 1065
rect -9725 1050 -9675 1065
rect -9635 1050 -9585 1065
rect -9545 1050 -9495 1065
rect -9455 1050 -9405 1065
rect -9365 1050 -9315 1065
rect -9275 1050 -9225 1065
rect -9185 1050 -9135 1065
rect -9095 1050 -9045 1065
rect -9005 1050 -8955 1065
rect -8915 1050 -8865 1065
rect -8825 1050 -8775 1065
rect -8735 1050 -8685 1065
rect -8645 1050 -8595 1065
rect -8555 1050 -8505 1065
rect -8465 1050 -8415 1065
rect -8375 1050 -8325 1065
rect -8285 1050 -8235 1065
rect -8195 1050 -8145 1065
rect -8105 1050 -8055 1065
rect -8015 1050 -7965 1065
rect -7925 1050 -7875 1065
rect -7835 1050 -7785 1065
rect -7745 1050 -7695 1065
rect -7655 1050 -7605 1065
rect -7565 1050 -7515 1065
rect -7475 1050 -7425 1065
rect -7385 1050 -7335 1065
rect -7295 1050 -7245 1065
rect -7205 1050 -7155 1065
rect -7115 1050 -7065 1065
rect -7025 1050 -6975 1065
rect -6935 1050 -6885 1065
rect -6845 1050 -6795 1065
rect -6755 1050 -6705 1065
rect -6665 1050 -6615 1065
rect -6575 1050 -6525 1065
rect -6485 1050 -6435 1065
rect -6395 1050 -6345 1065
rect -6305 1050 -6255 1065
rect -6215 1050 -6165 1065
rect -6125 1050 -6075 1065
rect -6035 1050 -5985 1065
rect -5945 1050 -5895 1065
rect -5855 1050 -5805 1065
rect -5765 1050 -5715 1065
rect -5675 1050 -5625 1065
rect -5585 1050 -5535 1065
rect -5495 1050 -5445 1065
rect -5405 1050 -5355 1065
rect -5315 1050 -5265 1065
rect -5225 1050 -5175 1065
rect -5135 1050 -5085 1065
rect -5045 1050 -4995 1065
rect -4955 1050 -4905 1065
rect -4865 1050 -4815 1065
rect -4775 1050 -4725 1065
rect -4685 1050 -4635 1065
rect -4595 1050 -4545 1065
rect -4505 1050 -4455 1065
rect -4415 1050 -4365 1065
rect -4325 1050 -4275 1065
rect -4235 1050 -4185 1065
rect -4145 1050 -4095 1065
rect -4055 1050 -4005 1065
rect -3965 1050 -3915 1065
rect -3875 1050 -3825 1065
rect -3785 1050 -3735 1065
rect -3695 1050 -3645 1065
rect -3605 1050 -3555 1065
rect -3515 1050 -3465 1065
rect -3425 1050 -3375 1065
rect -3335 1050 -3285 1065
rect -3245 1050 -3195 1065
rect -3155 1050 -3105 1065
rect -3065 1050 -3015 1065
rect -2975 1050 -2925 1065
rect -2885 1050 -2835 1065
rect -2795 1050 -2745 1065
rect -2705 1050 -2655 1065
rect -2615 1050 -2565 1065
rect -2525 1050 -2475 1065
rect -2435 1050 -2385 1065
rect -2345 1050 -2295 1065
rect -2255 1050 -2205 1065
rect -2165 1050 -2115 1065
rect -2075 1050 -2025 1065
rect -1985 1050 -1935 1065
rect -1895 1050 -1845 1065
rect -1805 1050 -1755 1065
rect -1715 1050 -1665 1065
rect -1625 1050 -1575 1065
rect -1535 1050 -1485 1065
rect -1445 1050 -1395 1065
rect -1355 1050 -1305 1065
rect -1265 1050 -1215 1065
rect -1175 1050 -1125 1065
rect -1085 1050 -1035 1065
rect -995 1050 -945 1065
rect -905 1050 -855 1065
rect -815 1050 -765 1065
rect -725 1050 -675 1065
rect -635 1050 -585 1065
rect -545 1050 -495 1065
rect -455 1050 -405 1065
rect -365 1050 -315 1065
rect -275 1050 -225 1065
rect -185 1050 -135 1065
rect -95 1050 -45 1065
rect -11525 930 -11475 945
rect -11435 930 -11385 945
rect -11345 930 -11295 945
rect -11255 930 -11205 945
rect -11165 930 -11115 945
rect -11075 930 -11025 945
rect -10985 930 -10935 945
rect -10895 930 -10845 945
rect -10805 930 -10755 945
rect -10715 930 -10665 945
rect -10625 930 -10575 945
rect -10535 930 -10485 945
rect -10445 930 -10395 945
rect -10355 930 -10305 945
rect -10265 930 -10215 945
rect -10175 930 -10125 945
rect -10085 930 -10035 945
rect -9995 930 -9945 945
rect -9905 930 -9855 945
rect -9815 930 -9765 945
rect -9725 930 -9675 945
rect -9635 930 -9585 945
rect -9545 930 -9495 945
rect -9455 930 -9405 945
rect -9365 930 -9315 945
rect -9275 930 -9225 945
rect -9185 930 -9135 945
rect -9095 930 -9045 945
rect -9005 930 -8955 945
rect -8915 930 -8865 945
rect -8825 930 -8775 945
rect -8735 930 -8685 945
rect -8645 930 -8595 945
rect -8555 930 -8505 945
rect -8465 930 -8415 945
rect -8375 930 -8325 945
rect -8285 930 -8235 945
rect -8195 930 -8145 945
rect -8105 930 -8055 945
rect -8015 930 -7965 945
rect -7925 930 -7875 945
rect -7835 930 -7785 945
rect -7745 930 -7695 945
rect -7655 930 -7605 945
rect -7565 930 -7515 945
rect -7475 930 -7425 945
rect -7385 930 -7335 945
rect -7295 930 -7245 945
rect -7205 930 -7155 945
rect -7115 930 -7065 945
rect -7025 930 -6975 945
rect -6935 930 -6885 945
rect -6845 930 -6795 945
rect -6755 930 -6705 945
rect -6665 930 -6615 945
rect -6575 930 -6525 945
rect -6485 930 -6435 945
rect -6395 930 -6345 945
rect -6305 930 -6255 945
rect -6215 930 -6165 945
rect -6125 930 -6075 945
rect -6035 930 -5985 945
rect -5945 930 -5895 945
rect -5855 930 -5805 945
rect -5765 930 -5715 945
rect -5675 930 -5625 945
rect -5585 930 -5535 945
rect -5495 930 -5445 945
rect -5405 930 -5355 945
rect -5315 930 -5265 945
rect -5225 930 -5175 945
rect -5135 930 -5085 945
rect -5045 930 -4995 945
rect -4955 930 -4905 945
rect -4865 930 -4815 945
rect -4775 930 -4725 945
rect -4685 930 -4635 945
rect -4595 930 -4545 945
rect -4505 930 -4455 945
rect -4415 930 -4365 945
rect -4325 930 -4275 945
rect -4235 930 -4185 945
rect -4145 930 -4095 945
rect -4055 930 -4005 945
rect -3965 930 -3915 945
rect -3875 930 -3825 945
rect -3785 930 -3735 945
rect -3695 930 -3645 945
rect -3605 930 -3555 945
rect -3515 930 -3465 945
rect -3425 930 -3375 945
rect -3335 930 -3285 945
rect -3245 930 -3195 945
rect -3155 930 -3105 945
rect -3065 930 -3015 945
rect -2975 930 -2925 945
rect -2885 930 -2835 945
rect -2795 930 -2745 945
rect -2705 930 -2655 945
rect -2615 930 -2565 945
rect -2525 930 -2475 945
rect -2435 930 -2385 945
rect -2345 930 -2295 945
rect -2255 930 -2205 945
rect -2165 930 -2115 945
rect -2075 930 -2025 945
rect -1985 930 -1935 945
rect -1895 930 -1845 945
rect -1805 930 -1755 945
rect -1715 930 -1665 945
rect -1625 930 -1575 945
rect -1535 930 -1485 945
rect -1445 930 -1395 945
rect -1355 930 -1305 945
rect -1265 930 -1215 945
rect -1175 930 -1125 945
rect -1085 930 -1035 945
rect -995 930 -945 945
rect -905 930 -855 945
rect -815 930 -765 945
rect -725 930 -675 945
rect -635 930 -585 945
rect -545 930 -495 945
rect -455 930 -405 945
rect -365 930 -315 945
rect -275 930 -225 945
rect -185 930 -135 945
rect -95 930 -45 945
rect -11525 810 -11475 830
rect -11435 810 -11385 830
rect -11525 805 -11385 810
rect -11525 785 -11510 805
rect -11490 785 -11420 805
rect -11400 785 -11385 805
rect -11525 780 -11385 785
rect -11345 810 -11295 830
rect -11255 810 -11205 830
rect -11345 805 -11205 810
rect -11345 785 -11330 805
rect -11310 785 -11240 805
rect -11220 785 -11205 805
rect -11345 780 -11205 785
rect -11165 810 -11115 830
rect -11075 810 -11025 830
rect -11165 805 -11025 810
rect -11165 785 -11150 805
rect -11130 785 -11060 805
rect -11040 785 -11025 805
rect -11165 780 -11025 785
rect -10985 810 -10935 830
rect -10895 810 -10845 830
rect -10985 805 -10845 810
rect -10985 785 -10970 805
rect -10950 785 -10880 805
rect -10860 785 -10845 805
rect -10985 780 -10845 785
rect -10805 810 -10755 830
rect -10715 810 -10665 830
rect -10805 805 -10665 810
rect -10805 785 -10790 805
rect -10770 785 -10700 805
rect -10680 785 -10665 805
rect -10805 780 -10665 785
rect -10625 810 -10575 830
rect -10535 810 -10485 830
rect -10625 805 -10485 810
rect -10625 785 -10610 805
rect -10590 785 -10520 805
rect -10500 785 -10485 805
rect -10625 780 -10485 785
rect -10445 810 -10395 830
rect -10355 810 -10305 830
rect -10445 805 -10305 810
rect -10445 785 -10430 805
rect -10410 785 -10340 805
rect -10320 785 -10305 805
rect -10445 780 -10305 785
rect -10265 810 -10215 830
rect -10175 810 -10125 830
rect -10265 805 -10125 810
rect -10265 785 -10250 805
rect -10230 785 -10160 805
rect -10140 785 -10125 805
rect -10265 780 -10125 785
rect -10085 810 -10035 830
rect -9995 810 -9945 830
rect -10085 805 -9945 810
rect -10085 785 -10070 805
rect -10050 785 -9980 805
rect -9960 785 -9945 805
rect -10085 780 -9945 785
rect -9905 810 -9855 830
rect -9815 810 -9765 830
rect -9905 805 -9765 810
rect -9905 785 -9890 805
rect -9870 785 -9800 805
rect -9780 785 -9765 805
rect -9905 780 -9765 785
rect -9725 810 -9675 830
rect -9635 810 -9585 830
rect -9725 805 -9585 810
rect -9725 785 -9710 805
rect -9690 785 -9620 805
rect -9600 785 -9585 805
rect -9725 780 -9585 785
rect -9545 810 -9495 830
rect -9455 810 -9405 830
rect -9545 805 -9405 810
rect -9545 785 -9530 805
rect -9510 785 -9440 805
rect -9420 785 -9405 805
rect -9545 780 -9405 785
rect -9365 810 -9315 830
rect -9275 810 -9225 830
rect -9365 805 -9225 810
rect -9365 785 -9350 805
rect -9330 785 -9260 805
rect -9240 785 -9225 805
rect -9365 780 -9225 785
rect -9185 810 -9135 830
rect -9095 810 -9045 830
rect -9185 805 -9045 810
rect -9185 785 -9170 805
rect -9150 785 -9080 805
rect -9060 785 -9045 805
rect -9185 780 -9045 785
rect -9005 810 -8955 830
rect -8915 810 -8865 830
rect -9005 805 -8865 810
rect -9005 785 -8990 805
rect -8970 785 -8900 805
rect -8880 785 -8865 805
rect -9005 780 -8865 785
rect -8825 810 -8775 830
rect -8735 810 -8685 830
rect -8825 805 -8685 810
rect -8825 785 -8810 805
rect -8790 785 -8720 805
rect -8700 785 -8685 805
rect -8825 780 -8685 785
rect -8645 810 -8595 830
rect -8555 810 -8505 830
rect -8645 805 -8505 810
rect -8645 785 -8630 805
rect -8610 785 -8540 805
rect -8520 785 -8505 805
rect -8645 780 -8505 785
rect -8465 810 -8415 830
rect -8375 810 -8325 830
rect -8465 805 -8325 810
rect -8465 785 -8450 805
rect -8430 785 -8360 805
rect -8340 785 -8325 805
rect -8465 780 -8325 785
rect -8285 810 -8235 830
rect -8195 810 -8145 830
rect -8285 805 -8145 810
rect -8285 785 -8270 805
rect -8250 785 -8180 805
rect -8160 785 -8145 805
rect -8285 780 -8145 785
rect -8105 810 -8055 830
rect -8015 810 -7965 830
rect -8105 805 -7965 810
rect -8105 785 -8090 805
rect -8070 785 -8000 805
rect -7980 785 -7965 805
rect -8105 780 -7965 785
rect -7925 810 -7875 830
rect -7835 810 -7785 830
rect -7925 805 -7785 810
rect -7925 785 -7910 805
rect -7890 785 -7820 805
rect -7800 785 -7785 805
rect -7925 780 -7785 785
rect -7745 810 -7695 830
rect -7655 810 -7605 830
rect -7745 805 -7605 810
rect -7745 785 -7730 805
rect -7710 785 -7640 805
rect -7620 785 -7605 805
rect -7745 780 -7605 785
rect -7565 810 -7515 830
rect -7475 810 -7425 830
rect -7565 805 -7425 810
rect -7565 785 -7550 805
rect -7530 785 -7460 805
rect -7440 785 -7425 805
rect -7565 780 -7425 785
rect -7385 810 -7335 830
rect -7295 810 -7245 830
rect -7385 805 -7245 810
rect -7385 785 -7370 805
rect -7350 785 -7280 805
rect -7260 785 -7245 805
rect -7385 780 -7245 785
rect -7205 810 -7155 830
rect -7115 810 -7065 830
rect -7205 805 -7065 810
rect -7205 785 -7190 805
rect -7170 785 -7100 805
rect -7080 785 -7065 805
rect -7205 780 -7065 785
rect -7025 810 -6975 830
rect -6935 810 -6885 830
rect -7025 805 -6885 810
rect -7025 785 -7010 805
rect -6990 785 -6920 805
rect -6900 785 -6885 805
rect -7025 780 -6885 785
rect -6845 810 -6795 830
rect -6755 810 -6705 830
rect -6845 805 -6705 810
rect -6845 785 -6830 805
rect -6810 785 -6740 805
rect -6720 785 -6705 805
rect -6845 780 -6705 785
rect -6665 810 -6615 830
rect -6575 810 -6525 830
rect -6665 805 -6525 810
rect -6665 785 -6650 805
rect -6630 785 -6560 805
rect -6540 785 -6525 805
rect -6665 780 -6525 785
rect -6485 810 -6435 830
rect -6395 810 -6345 830
rect -6485 805 -6345 810
rect -6485 785 -6470 805
rect -6450 785 -6380 805
rect -6360 785 -6345 805
rect -6485 780 -6345 785
rect -6305 810 -6255 830
rect -6215 810 -6165 830
rect -6305 805 -6165 810
rect -6305 785 -6290 805
rect -6270 785 -6200 805
rect -6180 785 -6165 805
rect -6305 780 -6165 785
rect -6125 810 -6075 830
rect -6035 810 -5985 830
rect -6125 805 -5985 810
rect -6125 785 -6110 805
rect -6090 785 -6020 805
rect -6000 785 -5985 805
rect -6125 780 -5985 785
rect -5945 810 -5895 830
rect -5855 810 -5805 830
rect -5945 805 -5805 810
rect -5945 785 -5930 805
rect -5910 785 -5840 805
rect -5820 785 -5805 805
rect -5945 780 -5805 785
rect -5765 810 -5715 830
rect -5675 810 -5625 830
rect -5765 805 -5625 810
rect -5765 785 -5750 805
rect -5730 785 -5660 805
rect -5640 785 -5625 805
rect -5765 780 -5625 785
rect -5585 810 -5535 830
rect -5495 810 -5445 830
rect -5585 805 -5445 810
rect -5585 785 -5570 805
rect -5550 785 -5480 805
rect -5460 785 -5445 805
rect -5585 780 -5445 785
rect -5405 810 -5355 830
rect -5315 810 -5265 830
rect -5405 805 -5265 810
rect -5405 785 -5390 805
rect -5370 785 -5300 805
rect -5280 785 -5265 805
rect -5405 780 -5265 785
rect -5225 810 -5175 830
rect -5135 810 -5085 830
rect -5225 805 -5085 810
rect -5225 785 -5210 805
rect -5190 785 -5120 805
rect -5100 785 -5085 805
rect -5225 780 -5085 785
rect -5045 810 -4995 830
rect -4955 810 -4905 830
rect -5045 805 -4905 810
rect -5045 785 -5030 805
rect -5010 785 -4940 805
rect -4920 785 -4905 805
rect -5045 780 -4905 785
rect -4865 810 -4815 830
rect -4775 810 -4725 830
rect -4865 805 -4725 810
rect -4865 785 -4850 805
rect -4830 785 -4760 805
rect -4740 785 -4725 805
rect -4865 780 -4725 785
rect -4685 810 -4635 830
rect -4595 810 -4545 830
rect -4685 805 -4545 810
rect -4685 785 -4670 805
rect -4650 785 -4580 805
rect -4560 785 -4545 805
rect -4685 780 -4545 785
rect -4505 810 -4455 830
rect -4415 810 -4365 830
rect -4505 805 -4365 810
rect -4505 785 -4490 805
rect -4470 785 -4400 805
rect -4380 785 -4365 805
rect -4505 780 -4365 785
rect -4325 810 -4275 830
rect -4235 810 -4185 830
rect -4325 805 -4185 810
rect -4325 785 -4310 805
rect -4290 785 -4220 805
rect -4200 785 -4185 805
rect -4325 780 -4185 785
rect -4145 810 -4095 830
rect -4055 810 -4005 830
rect -4145 805 -4005 810
rect -4145 785 -4130 805
rect -4110 785 -4040 805
rect -4020 785 -4005 805
rect -4145 780 -4005 785
rect -3965 810 -3915 830
rect -3875 810 -3825 830
rect -3965 805 -3825 810
rect -3965 785 -3950 805
rect -3930 785 -3860 805
rect -3840 785 -3825 805
rect -3965 780 -3825 785
rect -3785 810 -3735 830
rect -3695 810 -3645 830
rect -3785 805 -3645 810
rect -3785 785 -3770 805
rect -3750 785 -3680 805
rect -3660 785 -3645 805
rect -3785 780 -3645 785
rect -3605 810 -3555 830
rect -3515 810 -3465 830
rect -3605 805 -3465 810
rect -3605 785 -3590 805
rect -3570 785 -3500 805
rect -3480 785 -3465 805
rect -3605 780 -3465 785
rect -3425 810 -3375 830
rect -3335 810 -3285 830
rect -3425 805 -3285 810
rect -3425 785 -3410 805
rect -3390 785 -3320 805
rect -3300 785 -3285 805
rect -3425 780 -3285 785
rect -3245 810 -3195 830
rect -3155 810 -3105 830
rect -3245 805 -3105 810
rect -3245 785 -3230 805
rect -3210 785 -3140 805
rect -3120 785 -3105 805
rect -3245 780 -3105 785
rect -3065 810 -3015 830
rect -2975 810 -2925 830
rect -3065 805 -2925 810
rect -3065 785 -3050 805
rect -3030 785 -2960 805
rect -2940 785 -2925 805
rect -3065 780 -2925 785
rect -2885 810 -2835 830
rect -2795 810 -2745 830
rect -2885 805 -2745 810
rect -2885 785 -2870 805
rect -2850 785 -2780 805
rect -2760 785 -2745 805
rect -2885 780 -2745 785
rect -2705 810 -2655 830
rect -2615 810 -2565 830
rect -2705 805 -2565 810
rect -2705 785 -2690 805
rect -2670 785 -2600 805
rect -2580 785 -2565 805
rect -2705 780 -2565 785
rect -2525 810 -2475 830
rect -2435 810 -2385 830
rect -2525 805 -2385 810
rect -2525 785 -2510 805
rect -2490 785 -2420 805
rect -2400 785 -2385 805
rect -2525 780 -2385 785
rect -2345 810 -2295 830
rect -2255 810 -2205 830
rect -2345 805 -2205 810
rect -2345 785 -2330 805
rect -2310 785 -2240 805
rect -2220 785 -2205 805
rect -2345 780 -2205 785
rect -2165 810 -2115 830
rect -2075 810 -2025 830
rect -2165 805 -2025 810
rect -2165 785 -2150 805
rect -2130 785 -2060 805
rect -2040 785 -2025 805
rect -2165 780 -2025 785
rect -1985 810 -1935 830
rect -1895 810 -1845 830
rect -1985 805 -1845 810
rect -1985 785 -1970 805
rect -1950 785 -1880 805
rect -1860 785 -1845 805
rect -1985 780 -1845 785
rect -1805 810 -1755 830
rect -1715 810 -1665 830
rect -1805 805 -1665 810
rect -1805 785 -1790 805
rect -1770 785 -1700 805
rect -1680 785 -1665 805
rect -1805 780 -1665 785
rect -1625 810 -1575 830
rect -1535 810 -1485 830
rect -1625 805 -1485 810
rect -1625 785 -1610 805
rect -1590 785 -1520 805
rect -1500 785 -1485 805
rect -1625 780 -1485 785
rect -1445 810 -1395 830
rect -1355 810 -1305 830
rect -1445 805 -1305 810
rect -1445 785 -1430 805
rect -1410 785 -1340 805
rect -1320 785 -1305 805
rect -1445 780 -1305 785
rect -1265 810 -1215 830
rect -1175 810 -1125 830
rect -1265 805 -1125 810
rect -1265 785 -1250 805
rect -1230 785 -1160 805
rect -1140 785 -1125 805
rect -1265 780 -1125 785
rect -1085 810 -1035 830
rect -995 810 -945 830
rect -1085 805 -945 810
rect -1085 785 -1070 805
rect -1050 785 -980 805
rect -960 785 -945 805
rect -1085 780 -945 785
rect -905 810 -855 830
rect -815 810 -765 830
rect -905 805 -765 810
rect -905 785 -890 805
rect -870 785 -800 805
rect -780 785 -765 805
rect -905 780 -765 785
rect -725 810 -675 830
rect -635 810 -585 830
rect -725 805 -585 810
rect -725 785 -710 805
rect -690 785 -620 805
rect -600 785 -585 805
rect -725 780 -585 785
rect -545 810 -495 830
rect -455 810 -405 830
rect -545 805 -405 810
rect -545 785 -530 805
rect -510 785 -440 805
rect -420 785 -405 805
rect -545 780 -405 785
rect -365 810 -315 830
rect -275 810 -225 830
rect -365 805 -225 810
rect -365 785 -350 805
rect -330 785 -260 805
rect -240 785 -225 805
rect -365 780 -225 785
rect -185 810 -135 830
rect -95 810 -45 830
rect -185 805 -45 810
rect -185 785 -170 805
rect -150 785 -80 805
rect -60 785 -45 805
rect -185 780 -45 785
rect -11525 195 -11385 200
rect -11525 175 -11510 195
rect -11490 175 -11420 195
rect -11400 175 -11385 195
rect -11525 170 -11385 175
rect -11525 150 -11475 170
rect -11435 150 -11385 170
rect -11345 195 -11205 200
rect -11345 175 -11330 195
rect -11310 175 -11240 195
rect -11220 175 -11205 195
rect -11345 170 -11205 175
rect -11345 150 -11295 170
rect -11255 150 -11205 170
rect -11165 195 -11025 200
rect -11165 175 -11150 195
rect -11130 175 -11060 195
rect -11040 175 -11025 195
rect -11165 170 -11025 175
rect -11165 150 -11115 170
rect -11075 150 -11025 170
rect -10985 195 -10845 200
rect -10985 175 -10970 195
rect -10950 175 -10880 195
rect -10860 175 -10845 195
rect -10985 170 -10845 175
rect -10985 150 -10935 170
rect -10895 150 -10845 170
rect -10805 195 -10665 200
rect -10805 175 -10790 195
rect -10770 175 -10700 195
rect -10680 175 -10665 195
rect -10805 170 -10665 175
rect -10805 150 -10755 170
rect -10715 150 -10665 170
rect -10625 195 -10485 200
rect -10625 175 -10610 195
rect -10590 175 -10520 195
rect -10500 175 -10485 195
rect -10625 170 -10485 175
rect -10625 150 -10575 170
rect -10535 150 -10485 170
rect -10445 195 -10305 200
rect -10445 175 -10430 195
rect -10410 175 -10340 195
rect -10320 175 -10305 195
rect -10445 170 -10305 175
rect -10445 150 -10395 170
rect -10355 150 -10305 170
rect -10265 195 -10125 200
rect -10265 175 -10250 195
rect -10230 175 -10160 195
rect -10140 175 -10125 195
rect -10265 170 -10125 175
rect -10265 150 -10215 170
rect -10175 150 -10125 170
rect -10085 195 -9945 200
rect -10085 175 -10070 195
rect -10050 175 -9980 195
rect -9960 175 -9945 195
rect -10085 170 -9945 175
rect -10085 150 -10035 170
rect -9995 150 -9945 170
rect -9905 195 -9765 200
rect -9905 175 -9890 195
rect -9870 175 -9800 195
rect -9780 175 -9765 195
rect -9905 170 -9765 175
rect -9905 150 -9855 170
rect -9815 150 -9765 170
rect -9725 195 -9585 200
rect -9725 175 -9710 195
rect -9690 175 -9620 195
rect -9600 175 -9585 195
rect -9725 170 -9585 175
rect -9725 150 -9675 170
rect -9635 150 -9585 170
rect -9545 195 -9405 200
rect -9545 175 -9530 195
rect -9510 175 -9440 195
rect -9420 175 -9405 195
rect -9545 170 -9405 175
rect -9545 150 -9495 170
rect -9455 150 -9405 170
rect -9365 195 -9225 200
rect -9365 175 -9350 195
rect -9330 175 -9260 195
rect -9240 175 -9225 195
rect -9365 170 -9225 175
rect -9365 150 -9315 170
rect -9275 150 -9225 170
rect -9185 195 -9045 200
rect -9185 175 -9170 195
rect -9150 175 -9080 195
rect -9060 175 -9045 195
rect -9185 170 -9045 175
rect -9185 150 -9135 170
rect -9095 150 -9045 170
rect -9005 195 -8865 200
rect -9005 175 -8990 195
rect -8970 175 -8900 195
rect -8880 175 -8865 195
rect -9005 170 -8865 175
rect -9005 150 -8955 170
rect -8915 150 -8865 170
rect -8825 195 -8685 200
rect -8825 175 -8810 195
rect -8790 175 -8720 195
rect -8700 175 -8685 195
rect -8825 170 -8685 175
rect -8825 150 -8775 170
rect -8735 150 -8685 170
rect -8645 195 -8505 200
rect -8645 175 -8630 195
rect -8610 175 -8540 195
rect -8520 175 -8505 195
rect -8645 170 -8505 175
rect -8645 150 -8595 170
rect -8555 150 -8505 170
rect -8465 195 -8325 200
rect -8465 175 -8450 195
rect -8430 175 -8360 195
rect -8340 175 -8325 195
rect -8465 170 -8325 175
rect -8465 150 -8415 170
rect -8375 150 -8325 170
rect -8285 195 -8145 200
rect -8285 175 -8270 195
rect -8250 175 -8180 195
rect -8160 175 -8145 195
rect -8285 170 -8145 175
rect -8285 150 -8235 170
rect -8195 150 -8145 170
rect -8105 195 -7965 200
rect -8105 175 -8090 195
rect -8070 175 -8000 195
rect -7980 175 -7965 195
rect -8105 170 -7965 175
rect -8105 150 -8055 170
rect -8015 150 -7965 170
rect -7925 195 -7785 200
rect -7925 175 -7910 195
rect -7890 175 -7820 195
rect -7800 175 -7785 195
rect -7925 170 -7785 175
rect -7925 150 -7875 170
rect -7835 150 -7785 170
rect -7745 195 -7605 200
rect -7745 175 -7730 195
rect -7710 175 -7640 195
rect -7620 175 -7605 195
rect -7745 170 -7605 175
rect -7745 150 -7695 170
rect -7655 150 -7605 170
rect -7565 195 -7425 200
rect -7565 175 -7550 195
rect -7530 175 -7460 195
rect -7440 175 -7425 195
rect -7565 170 -7425 175
rect -7565 150 -7515 170
rect -7475 150 -7425 170
rect -7385 195 -7245 200
rect -7385 175 -7370 195
rect -7350 175 -7280 195
rect -7260 175 -7245 195
rect -7385 170 -7245 175
rect -7385 150 -7335 170
rect -7295 150 -7245 170
rect -7205 195 -7065 200
rect -7205 175 -7190 195
rect -7170 175 -7100 195
rect -7080 175 -7065 195
rect -7205 170 -7065 175
rect -7205 150 -7155 170
rect -7115 150 -7065 170
rect -7025 195 -6885 200
rect -7025 175 -7010 195
rect -6990 175 -6920 195
rect -6900 175 -6885 195
rect -7025 170 -6885 175
rect -7025 150 -6975 170
rect -6935 150 -6885 170
rect -6845 195 -6705 200
rect -6845 175 -6830 195
rect -6810 175 -6740 195
rect -6720 175 -6705 195
rect -6845 170 -6705 175
rect -6845 150 -6795 170
rect -6755 150 -6705 170
rect -6665 195 -6525 200
rect -6665 175 -6650 195
rect -6630 175 -6560 195
rect -6540 175 -6525 195
rect -6665 170 -6525 175
rect -6665 150 -6615 170
rect -6575 150 -6525 170
rect -6485 195 -6345 200
rect -6485 175 -6470 195
rect -6450 175 -6380 195
rect -6360 175 -6345 195
rect -6485 170 -6345 175
rect -6485 150 -6435 170
rect -6395 150 -6345 170
rect -6305 195 -6165 200
rect -6305 175 -6290 195
rect -6270 175 -6200 195
rect -6180 175 -6165 195
rect -6305 170 -6165 175
rect -6305 150 -6255 170
rect -6215 150 -6165 170
rect -6125 195 -5985 200
rect -6125 175 -6110 195
rect -6090 175 -6020 195
rect -6000 175 -5985 195
rect -6125 170 -5985 175
rect -6125 150 -6075 170
rect -6035 150 -5985 170
rect -5945 195 -5805 200
rect -5945 175 -5930 195
rect -5910 175 -5840 195
rect -5820 175 -5805 195
rect -5945 170 -5805 175
rect -5945 150 -5895 170
rect -5855 150 -5805 170
rect -5765 195 -5625 200
rect -5765 175 -5750 195
rect -5730 175 -5660 195
rect -5640 175 -5625 195
rect -5765 170 -5625 175
rect -5765 150 -5715 170
rect -5675 150 -5625 170
rect -5585 195 -5445 200
rect -5585 175 -5570 195
rect -5550 175 -5480 195
rect -5460 175 -5445 195
rect -5585 170 -5445 175
rect -5585 150 -5535 170
rect -5495 150 -5445 170
rect -5405 195 -5265 200
rect -5405 175 -5390 195
rect -5370 175 -5300 195
rect -5280 175 -5265 195
rect -5405 170 -5265 175
rect -5405 150 -5355 170
rect -5315 150 -5265 170
rect -5225 195 -5085 200
rect -5225 175 -5210 195
rect -5190 175 -5120 195
rect -5100 175 -5085 195
rect -5225 170 -5085 175
rect -5225 150 -5175 170
rect -5135 150 -5085 170
rect -5045 195 -4905 200
rect -5045 175 -5030 195
rect -5010 175 -4940 195
rect -4920 175 -4905 195
rect -5045 170 -4905 175
rect -5045 150 -4995 170
rect -4955 150 -4905 170
rect -4865 195 -4725 200
rect -4865 175 -4850 195
rect -4830 175 -4760 195
rect -4740 175 -4725 195
rect -4865 170 -4725 175
rect -4865 150 -4815 170
rect -4775 150 -4725 170
rect -4685 195 -4545 200
rect -4685 175 -4670 195
rect -4650 175 -4580 195
rect -4560 175 -4545 195
rect -4685 170 -4545 175
rect -4685 150 -4635 170
rect -4595 150 -4545 170
rect -4505 195 -4365 200
rect -4505 175 -4490 195
rect -4470 175 -4400 195
rect -4380 175 -4365 195
rect -4505 170 -4365 175
rect -4505 150 -4455 170
rect -4415 150 -4365 170
rect -4325 195 -4185 200
rect -4325 175 -4310 195
rect -4290 175 -4220 195
rect -4200 175 -4185 195
rect -4325 170 -4185 175
rect -4325 150 -4275 170
rect -4235 150 -4185 170
rect -4145 195 -4005 200
rect -4145 175 -4130 195
rect -4110 175 -4040 195
rect -4020 175 -4005 195
rect -4145 170 -4005 175
rect -4145 150 -4095 170
rect -4055 150 -4005 170
rect -3965 195 -3825 200
rect -3965 175 -3950 195
rect -3930 175 -3860 195
rect -3840 175 -3825 195
rect -3965 170 -3825 175
rect -3965 150 -3915 170
rect -3875 150 -3825 170
rect -3785 195 -3645 200
rect -3785 175 -3770 195
rect -3750 175 -3680 195
rect -3660 175 -3645 195
rect -3785 170 -3645 175
rect -3785 150 -3735 170
rect -3695 150 -3645 170
rect -3605 195 -3465 200
rect -3605 175 -3590 195
rect -3570 175 -3500 195
rect -3480 175 -3465 195
rect -3605 170 -3465 175
rect -3605 150 -3555 170
rect -3515 150 -3465 170
rect -3425 195 -3285 200
rect -3425 175 -3410 195
rect -3390 175 -3320 195
rect -3300 175 -3285 195
rect -3425 170 -3285 175
rect -3425 150 -3375 170
rect -3335 150 -3285 170
rect -3245 195 -3105 200
rect -3245 175 -3230 195
rect -3210 175 -3140 195
rect -3120 175 -3105 195
rect -3245 170 -3105 175
rect -3245 150 -3195 170
rect -3155 150 -3105 170
rect -3065 195 -2925 200
rect -3065 175 -3050 195
rect -3030 175 -2960 195
rect -2940 175 -2925 195
rect -3065 170 -2925 175
rect -3065 150 -3015 170
rect -2975 150 -2925 170
rect -2885 195 -2745 200
rect -2885 175 -2870 195
rect -2850 175 -2780 195
rect -2760 175 -2745 195
rect -2885 170 -2745 175
rect -2885 150 -2835 170
rect -2795 150 -2745 170
rect -2705 195 -2565 200
rect -2705 175 -2690 195
rect -2670 175 -2600 195
rect -2580 175 -2565 195
rect -2705 170 -2565 175
rect -2705 150 -2655 170
rect -2615 150 -2565 170
rect -2525 195 -2385 200
rect -2525 175 -2510 195
rect -2490 175 -2420 195
rect -2400 175 -2385 195
rect -2525 170 -2385 175
rect -2525 150 -2475 170
rect -2435 150 -2385 170
rect -2345 195 -2205 200
rect -2345 175 -2330 195
rect -2310 175 -2240 195
rect -2220 175 -2205 195
rect -2345 170 -2205 175
rect -2345 150 -2295 170
rect -2255 150 -2205 170
rect -2165 195 -2025 200
rect -2165 175 -2150 195
rect -2130 175 -2060 195
rect -2040 175 -2025 195
rect -2165 170 -2025 175
rect -2165 150 -2115 170
rect -2075 150 -2025 170
rect -1985 195 -1845 200
rect -1985 175 -1970 195
rect -1950 175 -1880 195
rect -1860 175 -1845 195
rect -1985 170 -1845 175
rect -1985 150 -1935 170
rect -1895 150 -1845 170
rect -1805 195 -1665 200
rect -1805 175 -1790 195
rect -1770 175 -1700 195
rect -1680 175 -1665 195
rect -1805 170 -1665 175
rect -1805 150 -1755 170
rect -1715 150 -1665 170
rect -1625 195 -1485 200
rect -1625 175 -1610 195
rect -1590 175 -1520 195
rect -1500 175 -1485 195
rect -1625 170 -1485 175
rect -1625 150 -1575 170
rect -1535 150 -1485 170
rect -1445 195 -1305 200
rect -1445 175 -1430 195
rect -1410 175 -1340 195
rect -1320 175 -1305 195
rect -1445 170 -1305 175
rect -1445 150 -1395 170
rect -1355 150 -1305 170
rect -1265 195 -1125 200
rect -1265 175 -1250 195
rect -1230 175 -1160 195
rect -1140 175 -1125 195
rect -1265 170 -1125 175
rect -1265 150 -1215 170
rect -1175 150 -1125 170
rect -1085 195 -945 200
rect -1085 175 -1070 195
rect -1050 175 -980 195
rect -960 175 -945 195
rect -1085 170 -945 175
rect -1085 150 -1035 170
rect -995 150 -945 170
rect -905 195 -765 200
rect -905 175 -890 195
rect -870 175 -800 195
rect -780 175 -765 195
rect -905 170 -765 175
rect -905 150 -855 170
rect -815 150 -765 170
rect -725 195 -585 200
rect -725 175 -710 195
rect -690 175 -620 195
rect -600 175 -585 195
rect -725 170 -585 175
rect -725 150 -675 170
rect -635 150 -585 170
rect -545 195 -405 200
rect -545 175 -530 195
rect -510 175 -440 195
rect -420 175 -405 195
rect -545 170 -405 175
rect -545 150 -495 170
rect -455 150 -405 170
rect -365 195 -225 200
rect -365 175 -350 195
rect -330 175 -260 195
rect -240 175 -225 195
rect -365 170 -225 175
rect -365 150 -315 170
rect -275 150 -225 170
rect -185 195 -45 200
rect -185 175 -170 195
rect -150 175 -80 195
rect -60 175 -45 195
rect -185 170 -45 175
rect -185 150 -135 170
rect -95 150 -45 170
rect -11525 35 -11475 50
rect -11435 35 -11385 50
rect -11345 35 -11295 50
rect -11255 35 -11205 50
rect -11165 35 -11115 50
rect -11075 35 -11025 50
rect -10985 35 -10935 50
rect -10895 35 -10845 50
rect -10805 35 -10755 50
rect -10715 35 -10665 50
rect -10625 35 -10575 50
rect -10535 35 -10485 50
rect -10445 35 -10395 50
rect -10355 35 -10305 50
rect -10265 35 -10215 50
rect -10175 35 -10125 50
rect -10085 35 -10035 50
rect -9995 35 -9945 50
rect -9905 35 -9855 50
rect -9815 35 -9765 50
rect -9725 35 -9675 50
rect -9635 35 -9585 50
rect -9545 35 -9495 50
rect -9455 35 -9405 50
rect -9365 35 -9315 50
rect -9275 35 -9225 50
rect -9185 35 -9135 50
rect -9095 35 -9045 50
rect -9005 35 -8955 50
rect -8915 35 -8865 50
rect -8825 35 -8775 50
rect -8735 35 -8685 50
rect -8645 35 -8595 50
rect -8555 35 -8505 50
rect -8465 35 -8415 50
rect -8375 35 -8325 50
rect -8285 35 -8235 50
rect -8195 35 -8145 50
rect -8105 35 -8055 50
rect -8015 35 -7965 50
rect -7925 35 -7875 50
rect -7835 35 -7785 50
rect -7745 35 -7695 50
rect -7655 35 -7605 50
rect -7565 35 -7515 50
rect -7475 35 -7425 50
rect -7385 35 -7335 50
rect -7295 35 -7245 50
rect -7205 35 -7155 50
rect -7115 35 -7065 50
rect -7025 35 -6975 50
rect -6935 35 -6885 50
rect -6845 35 -6795 50
rect -6755 35 -6705 50
rect -6665 35 -6615 50
rect -6575 35 -6525 50
rect -6485 35 -6435 50
rect -6395 35 -6345 50
rect -6305 35 -6255 50
rect -6215 35 -6165 50
rect -6125 35 -6075 50
rect -6035 35 -5985 50
rect -5945 35 -5895 50
rect -5855 35 -5805 50
rect -5765 35 -5715 50
rect -5675 35 -5625 50
rect -5585 35 -5535 50
rect -5495 35 -5445 50
rect -5405 35 -5355 50
rect -5315 35 -5265 50
rect -5225 35 -5175 50
rect -5135 35 -5085 50
rect -5045 35 -4995 50
rect -4955 35 -4905 50
rect -4865 35 -4815 50
rect -4775 35 -4725 50
rect -4685 35 -4635 50
rect -4595 35 -4545 50
rect -4505 35 -4455 50
rect -4415 35 -4365 50
rect -4325 35 -4275 50
rect -4235 35 -4185 50
rect -4145 35 -4095 50
rect -4055 35 -4005 50
rect -3965 35 -3915 50
rect -3875 35 -3825 50
rect -3785 35 -3735 50
rect -3695 35 -3645 50
rect -3605 35 -3555 50
rect -3515 35 -3465 50
rect -3425 35 -3375 50
rect -3335 35 -3285 50
rect -3245 35 -3195 50
rect -3155 35 -3105 50
rect -3065 35 -3015 50
rect -2975 35 -2925 50
rect -2885 35 -2835 50
rect -2795 35 -2745 50
rect -2705 35 -2655 50
rect -2615 35 -2565 50
rect -2525 35 -2475 50
rect -2435 35 -2385 50
rect -2345 35 -2295 50
rect -2255 35 -2205 50
rect -2165 35 -2115 50
rect -2075 35 -2025 50
rect -1985 35 -1935 50
rect -1895 35 -1845 50
rect -1805 35 -1755 50
rect -1715 35 -1665 50
rect -1625 35 -1575 50
rect -1535 35 -1485 50
rect -1445 35 -1395 50
rect -1355 35 -1305 50
rect -1265 35 -1215 50
rect -1175 35 -1125 50
rect -1085 35 -1035 50
rect -995 35 -945 50
rect -905 35 -855 50
rect -815 35 -765 50
rect -725 35 -675 50
rect -635 35 -585 50
rect -545 35 -495 50
rect -455 35 -405 50
rect -365 35 -315 50
rect -275 35 -225 50
rect -185 35 -135 50
rect -95 35 -45 50
<< polycont >>
rect -11510 1800 -11490 1820
rect -11420 1800 -11400 1820
rect -11330 1800 -11310 1820
rect -11240 1800 -11220 1820
rect -11150 1800 -11130 1820
rect -11060 1800 -11040 1820
rect -10970 1800 -10950 1820
rect -10880 1800 -10860 1820
rect -10790 1800 -10770 1820
rect -10700 1800 -10680 1820
rect -10610 1800 -10590 1820
rect -10520 1800 -10500 1820
rect -10430 1800 -10410 1820
rect -10340 1800 -10320 1820
rect -10250 1800 -10230 1820
rect -10160 1800 -10140 1820
rect -10070 1800 -10050 1820
rect -9980 1800 -9960 1820
rect -9890 1800 -9870 1820
rect -9800 1800 -9780 1820
rect -9710 1800 -9690 1820
rect -9620 1800 -9600 1820
rect -9530 1800 -9510 1820
rect -9440 1800 -9420 1820
rect -9350 1800 -9330 1820
rect -9260 1800 -9240 1820
rect -9170 1800 -9150 1820
rect -9080 1800 -9060 1820
rect -8990 1800 -8970 1820
rect -8900 1800 -8880 1820
rect -8810 1800 -8790 1820
rect -8720 1800 -8700 1820
rect -8630 1800 -8610 1820
rect -8540 1800 -8520 1820
rect -8450 1800 -8430 1820
rect -8360 1800 -8340 1820
rect -8270 1800 -8250 1820
rect -8180 1800 -8160 1820
rect -8090 1800 -8070 1820
rect -8000 1800 -7980 1820
rect -7910 1800 -7890 1820
rect -7820 1800 -7800 1820
rect -7730 1800 -7710 1820
rect -7640 1800 -7620 1820
rect -7550 1800 -7530 1820
rect -7460 1800 -7440 1820
rect -7370 1800 -7350 1820
rect -7280 1800 -7260 1820
rect -7190 1800 -7170 1820
rect -7100 1800 -7080 1820
rect -7010 1800 -6990 1820
rect -6920 1800 -6900 1820
rect -6830 1800 -6810 1820
rect -6740 1800 -6720 1820
rect -6650 1800 -6630 1820
rect -6560 1800 -6540 1820
rect -6470 1800 -6450 1820
rect -6380 1800 -6360 1820
rect -6290 1800 -6270 1820
rect -6200 1800 -6180 1820
rect -6110 1800 -6090 1820
rect -6020 1800 -6000 1820
rect -5930 1800 -5910 1820
rect -5840 1800 -5820 1820
rect -5750 1800 -5730 1820
rect -5660 1800 -5640 1820
rect -5570 1800 -5550 1820
rect -5480 1800 -5460 1820
rect -5390 1800 -5370 1820
rect -5300 1800 -5280 1820
rect -5210 1800 -5190 1820
rect -5120 1800 -5100 1820
rect -5030 1800 -5010 1820
rect -4940 1800 -4920 1820
rect -4850 1800 -4830 1820
rect -4760 1800 -4740 1820
rect -4670 1800 -4650 1820
rect -4580 1800 -4560 1820
rect -4490 1800 -4470 1820
rect -4400 1800 -4380 1820
rect -4310 1800 -4290 1820
rect -4220 1800 -4200 1820
rect -4130 1800 -4110 1820
rect -4040 1800 -4020 1820
rect -3950 1800 -3930 1820
rect -3860 1800 -3840 1820
rect -3770 1800 -3750 1820
rect -3680 1800 -3660 1820
rect -3590 1800 -3570 1820
rect -3500 1800 -3480 1820
rect -3410 1800 -3390 1820
rect -3320 1800 -3300 1820
rect -3230 1800 -3210 1820
rect -3140 1800 -3120 1820
rect -3050 1800 -3030 1820
rect -2960 1800 -2940 1820
rect -2870 1800 -2850 1820
rect -2780 1800 -2760 1820
rect -2690 1800 -2670 1820
rect -2600 1800 -2580 1820
rect -2510 1800 -2490 1820
rect -2420 1800 -2400 1820
rect -2330 1800 -2310 1820
rect -2240 1800 -2220 1820
rect -2150 1800 -2130 1820
rect -2060 1800 -2040 1820
rect -1970 1800 -1950 1820
rect -1880 1800 -1860 1820
rect -1790 1800 -1770 1820
rect -1700 1800 -1680 1820
rect -1610 1800 -1590 1820
rect -1520 1800 -1500 1820
rect -1430 1800 -1410 1820
rect -1340 1800 -1320 1820
rect -1250 1800 -1230 1820
rect -1160 1800 -1140 1820
rect -1070 1800 -1050 1820
rect -980 1800 -960 1820
rect -890 1800 -870 1820
rect -800 1800 -780 1820
rect -710 1800 -690 1820
rect -620 1800 -600 1820
rect -530 1800 -510 1820
rect -440 1800 -420 1820
rect -350 1800 -330 1820
rect -260 1800 -240 1820
rect -170 1800 -150 1820
rect -80 1800 -60 1820
rect -11510 1190 -11490 1210
rect -11420 1190 -11400 1210
rect -11330 1190 -11310 1210
rect -11240 1190 -11220 1210
rect -11150 1190 -11130 1210
rect -11060 1190 -11040 1210
rect -10970 1190 -10950 1210
rect -10880 1190 -10860 1210
rect -10790 1190 -10770 1210
rect -10700 1190 -10680 1210
rect -10610 1190 -10590 1210
rect -10520 1190 -10500 1210
rect -10430 1190 -10410 1210
rect -10340 1190 -10320 1210
rect -10250 1190 -10230 1210
rect -10160 1190 -10140 1210
rect -10070 1190 -10050 1210
rect -9980 1190 -9960 1210
rect -9890 1190 -9870 1210
rect -9800 1190 -9780 1210
rect -9710 1190 -9690 1210
rect -9620 1190 -9600 1210
rect -9530 1190 -9510 1210
rect -9440 1190 -9420 1210
rect -9350 1190 -9330 1210
rect -9260 1190 -9240 1210
rect -9170 1190 -9150 1210
rect -9080 1190 -9060 1210
rect -8990 1190 -8970 1210
rect -8900 1190 -8880 1210
rect -8810 1190 -8790 1210
rect -8720 1190 -8700 1210
rect -8630 1190 -8610 1210
rect -8540 1190 -8520 1210
rect -8450 1190 -8430 1210
rect -8360 1190 -8340 1210
rect -8270 1190 -8250 1210
rect -8180 1190 -8160 1210
rect -8090 1190 -8070 1210
rect -8000 1190 -7980 1210
rect -7910 1190 -7890 1210
rect -7820 1190 -7800 1210
rect -7730 1190 -7710 1210
rect -7640 1190 -7620 1210
rect -7550 1190 -7530 1210
rect -7460 1190 -7440 1210
rect -7370 1190 -7350 1210
rect -7280 1190 -7260 1210
rect -7190 1190 -7170 1210
rect -7100 1190 -7080 1210
rect -7010 1190 -6990 1210
rect -6920 1190 -6900 1210
rect -6830 1190 -6810 1210
rect -6740 1190 -6720 1210
rect -6650 1190 -6630 1210
rect -6560 1190 -6540 1210
rect -6470 1190 -6450 1210
rect -6380 1190 -6360 1210
rect -6290 1190 -6270 1210
rect -6200 1190 -6180 1210
rect -6110 1190 -6090 1210
rect -6020 1190 -6000 1210
rect -5930 1190 -5910 1210
rect -5840 1190 -5820 1210
rect -5750 1190 -5730 1210
rect -5660 1190 -5640 1210
rect -5570 1190 -5550 1210
rect -5480 1190 -5460 1210
rect -5390 1190 -5370 1210
rect -5300 1190 -5280 1210
rect -5210 1190 -5190 1210
rect -5120 1190 -5100 1210
rect -5030 1190 -5010 1210
rect -4940 1190 -4920 1210
rect -4850 1190 -4830 1210
rect -4760 1190 -4740 1210
rect -4670 1190 -4650 1210
rect -4580 1190 -4560 1210
rect -4490 1190 -4470 1210
rect -4400 1190 -4380 1210
rect -4310 1190 -4290 1210
rect -4220 1190 -4200 1210
rect -4130 1190 -4110 1210
rect -4040 1190 -4020 1210
rect -3950 1190 -3930 1210
rect -3860 1190 -3840 1210
rect -3770 1190 -3750 1210
rect -3680 1190 -3660 1210
rect -3590 1190 -3570 1210
rect -3500 1190 -3480 1210
rect -3410 1190 -3390 1210
rect -3320 1190 -3300 1210
rect -3230 1190 -3210 1210
rect -3140 1190 -3120 1210
rect -3050 1190 -3030 1210
rect -2960 1190 -2940 1210
rect -2870 1190 -2850 1210
rect -2780 1190 -2760 1210
rect -2690 1190 -2670 1210
rect -2600 1190 -2580 1210
rect -2510 1190 -2490 1210
rect -2420 1190 -2400 1210
rect -2330 1190 -2310 1210
rect -2240 1190 -2220 1210
rect -2150 1190 -2130 1210
rect -2060 1190 -2040 1210
rect -1970 1190 -1950 1210
rect -1880 1190 -1860 1210
rect -1790 1190 -1770 1210
rect -1700 1190 -1680 1210
rect -1610 1190 -1590 1210
rect -1520 1190 -1500 1210
rect -1430 1190 -1410 1210
rect -1340 1190 -1320 1210
rect -1250 1190 -1230 1210
rect -1160 1190 -1140 1210
rect -1070 1190 -1050 1210
rect -980 1190 -960 1210
rect -890 1190 -870 1210
rect -800 1190 -780 1210
rect -710 1190 -690 1210
rect -620 1190 -600 1210
rect -530 1190 -510 1210
rect -440 1190 -420 1210
rect -350 1190 -330 1210
rect -260 1190 -240 1210
rect -170 1190 -150 1210
rect -80 1190 -60 1210
rect -11510 785 -11490 805
rect -11420 785 -11400 805
rect -11330 785 -11310 805
rect -11240 785 -11220 805
rect -11150 785 -11130 805
rect -11060 785 -11040 805
rect -10970 785 -10950 805
rect -10880 785 -10860 805
rect -10790 785 -10770 805
rect -10700 785 -10680 805
rect -10610 785 -10590 805
rect -10520 785 -10500 805
rect -10430 785 -10410 805
rect -10340 785 -10320 805
rect -10250 785 -10230 805
rect -10160 785 -10140 805
rect -10070 785 -10050 805
rect -9980 785 -9960 805
rect -9890 785 -9870 805
rect -9800 785 -9780 805
rect -9710 785 -9690 805
rect -9620 785 -9600 805
rect -9530 785 -9510 805
rect -9440 785 -9420 805
rect -9350 785 -9330 805
rect -9260 785 -9240 805
rect -9170 785 -9150 805
rect -9080 785 -9060 805
rect -8990 785 -8970 805
rect -8900 785 -8880 805
rect -8810 785 -8790 805
rect -8720 785 -8700 805
rect -8630 785 -8610 805
rect -8540 785 -8520 805
rect -8450 785 -8430 805
rect -8360 785 -8340 805
rect -8270 785 -8250 805
rect -8180 785 -8160 805
rect -8090 785 -8070 805
rect -8000 785 -7980 805
rect -7910 785 -7890 805
rect -7820 785 -7800 805
rect -7730 785 -7710 805
rect -7640 785 -7620 805
rect -7550 785 -7530 805
rect -7460 785 -7440 805
rect -7370 785 -7350 805
rect -7280 785 -7260 805
rect -7190 785 -7170 805
rect -7100 785 -7080 805
rect -7010 785 -6990 805
rect -6920 785 -6900 805
rect -6830 785 -6810 805
rect -6740 785 -6720 805
rect -6650 785 -6630 805
rect -6560 785 -6540 805
rect -6470 785 -6450 805
rect -6380 785 -6360 805
rect -6290 785 -6270 805
rect -6200 785 -6180 805
rect -6110 785 -6090 805
rect -6020 785 -6000 805
rect -5930 785 -5910 805
rect -5840 785 -5820 805
rect -5750 785 -5730 805
rect -5660 785 -5640 805
rect -5570 785 -5550 805
rect -5480 785 -5460 805
rect -5390 785 -5370 805
rect -5300 785 -5280 805
rect -5210 785 -5190 805
rect -5120 785 -5100 805
rect -5030 785 -5010 805
rect -4940 785 -4920 805
rect -4850 785 -4830 805
rect -4760 785 -4740 805
rect -4670 785 -4650 805
rect -4580 785 -4560 805
rect -4490 785 -4470 805
rect -4400 785 -4380 805
rect -4310 785 -4290 805
rect -4220 785 -4200 805
rect -4130 785 -4110 805
rect -4040 785 -4020 805
rect -3950 785 -3930 805
rect -3860 785 -3840 805
rect -3770 785 -3750 805
rect -3680 785 -3660 805
rect -3590 785 -3570 805
rect -3500 785 -3480 805
rect -3410 785 -3390 805
rect -3320 785 -3300 805
rect -3230 785 -3210 805
rect -3140 785 -3120 805
rect -3050 785 -3030 805
rect -2960 785 -2940 805
rect -2870 785 -2850 805
rect -2780 785 -2760 805
rect -2690 785 -2670 805
rect -2600 785 -2580 805
rect -2510 785 -2490 805
rect -2420 785 -2400 805
rect -2330 785 -2310 805
rect -2240 785 -2220 805
rect -2150 785 -2130 805
rect -2060 785 -2040 805
rect -1970 785 -1950 805
rect -1880 785 -1860 805
rect -1790 785 -1770 805
rect -1700 785 -1680 805
rect -1610 785 -1590 805
rect -1520 785 -1500 805
rect -1430 785 -1410 805
rect -1340 785 -1320 805
rect -1250 785 -1230 805
rect -1160 785 -1140 805
rect -1070 785 -1050 805
rect -980 785 -960 805
rect -890 785 -870 805
rect -800 785 -780 805
rect -710 785 -690 805
rect -620 785 -600 805
rect -530 785 -510 805
rect -440 785 -420 805
rect -350 785 -330 805
rect -260 785 -240 805
rect -170 785 -150 805
rect -80 785 -60 805
rect -11510 175 -11490 195
rect -11420 175 -11400 195
rect -11330 175 -11310 195
rect -11240 175 -11220 195
rect -11150 175 -11130 195
rect -11060 175 -11040 195
rect -10970 175 -10950 195
rect -10880 175 -10860 195
rect -10790 175 -10770 195
rect -10700 175 -10680 195
rect -10610 175 -10590 195
rect -10520 175 -10500 195
rect -10430 175 -10410 195
rect -10340 175 -10320 195
rect -10250 175 -10230 195
rect -10160 175 -10140 195
rect -10070 175 -10050 195
rect -9980 175 -9960 195
rect -9890 175 -9870 195
rect -9800 175 -9780 195
rect -9710 175 -9690 195
rect -9620 175 -9600 195
rect -9530 175 -9510 195
rect -9440 175 -9420 195
rect -9350 175 -9330 195
rect -9260 175 -9240 195
rect -9170 175 -9150 195
rect -9080 175 -9060 195
rect -8990 175 -8970 195
rect -8900 175 -8880 195
rect -8810 175 -8790 195
rect -8720 175 -8700 195
rect -8630 175 -8610 195
rect -8540 175 -8520 195
rect -8450 175 -8430 195
rect -8360 175 -8340 195
rect -8270 175 -8250 195
rect -8180 175 -8160 195
rect -8090 175 -8070 195
rect -8000 175 -7980 195
rect -7910 175 -7890 195
rect -7820 175 -7800 195
rect -7730 175 -7710 195
rect -7640 175 -7620 195
rect -7550 175 -7530 195
rect -7460 175 -7440 195
rect -7370 175 -7350 195
rect -7280 175 -7260 195
rect -7190 175 -7170 195
rect -7100 175 -7080 195
rect -7010 175 -6990 195
rect -6920 175 -6900 195
rect -6830 175 -6810 195
rect -6740 175 -6720 195
rect -6650 175 -6630 195
rect -6560 175 -6540 195
rect -6470 175 -6450 195
rect -6380 175 -6360 195
rect -6290 175 -6270 195
rect -6200 175 -6180 195
rect -6110 175 -6090 195
rect -6020 175 -6000 195
rect -5930 175 -5910 195
rect -5840 175 -5820 195
rect -5750 175 -5730 195
rect -5660 175 -5640 195
rect -5570 175 -5550 195
rect -5480 175 -5460 195
rect -5390 175 -5370 195
rect -5300 175 -5280 195
rect -5210 175 -5190 195
rect -5120 175 -5100 195
rect -5030 175 -5010 195
rect -4940 175 -4920 195
rect -4850 175 -4830 195
rect -4760 175 -4740 195
rect -4670 175 -4650 195
rect -4580 175 -4560 195
rect -4490 175 -4470 195
rect -4400 175 -4380 195
rect -4310 175 -4290 195
rect -4220 175 -4200 195
rect -4130 175 -4110 195
rect -4040 175 -4020 195
rect -3950 175 -3930 195
rect -3860 175 -3840 195
rect -3770 175 -3750 195
rect -3680 175 -3660 195
rect -3590 175 -3570 195
rect -3500 175 -3480 195
rect -3410 175 -3390 195
rect -3320 175 -3300 195
rect -3230 175 -3210 195
rect -3140 175 -3120 195
rect -3050 175 -3030 195
rect -2960 175 -2940 195
rect -2870 175 -2850 195
rect -2780 175 -2760 195
rect -2690 175 -2670 195
rect -2600 175 -2580 195
rect -2510 175 -2490 195
rect -2420 175 -2400 195
rect -2330 175 -2310 195
rect -2240 175 -2220 195
rect -2150 175 -2130 195
rect -2060 175 -2040 195
rect -1970 175 -1950 195
rect -1880 175 -1860 195
rect -1790 175 -1770 195
rect -1700 175 -1680 195
rect -1610 175 -1590 195
rect -1520 175 -1500 195
rect -1430 175 -1410 195
rect -1340 175 -1320 195
rect -1250 175 -1230 195
rect -1160 175 -1140 195
rect -1070 175 -1050 195
rect -980 175 -960 195
rect -890 175 -870 195
rect -800 175 -780 195
rect -710 175 -690 195
rect -620 175 -600 195
rect -530 175 -510 195
rect -440 175 -420 195
rect -350 175 -330 195
rect -260 175 -240 195
rect -170 175 -150 195
rect -80 175 -60 195
<< locali >>
rect -11700 1975 -11690 1995
rect -11670 1975 -11555 1995
rect -11535 1975 -11510 1995
rect -11490 1975 -11420 1995
rect -11400 1975 -11330 1995
rect -11310 1975 -11240 1995
rect -11220 1975 -11150 1995
rect -11130 1975 -11060 1995
rect -11040 1975 -10970 1995
rect -10950 1975 -10880 1995
rect -10860 1975 -10835 1995
rect -10815 1975 -10790 1995
rect -10770 1975 -10700 1995
rect -10680 1975 -10655 1995
rect -10635 1975 -10610 1995
rect -10590 1975 -10520 1995
rect -10500 1975 -10475 1995
rect -10455 1975 -10430 1995
rect -10410 1975 -10340 1995
rect -10320 1975 -10295 1995
rect -10275 1975 -10250 1995
rect -10230 1975 -10160 1995
rect -10140 1975 -10115 1995
rect -10095 1975 -10070 1995
rect -10050 1975 -9980 1995
rect -9960 1975 -9935 1995
rect -9915 1975 -9890 1995
rect -9870 1975 -9800 1995
rect -9780 1975 -9755 1995
rect -9735 1975 -9710 1995
rect -9690 1975 -9620 1995
rect -9600 1975 -9575 1995
rect -9555 1975 -9530 1995
rect -9510 1975 -9440 1995
rect -9420 1975 -9395 1995
rect -9375 1975 -9350 1995
rect -9330 1975 -9260 1995
rect -9240 1975 -9215 1995
rect -9195 1975 -9170 1995
rect -9150 1975 -9080 1995
rect -9060 1975 -9035 1995
rect -9015 1975 -8990 1995
rect -8970 1975 -8900 1995
rect -8880 1975 -8855 1995
rect -8835 1975 -8810 1995
rect -8790 1975 -8720 1995
rect -8700 1975 -8675 1995
rect -8655 1975 -8630 1995
rect -8610 1975 -8540 1995
rect -8520 1975 -8495 1995
rect -8475 1975 -8450 1995
rect -8430 1975 -8360 1995
rect -8340 1975 -8315 1995
rect -8295 1975 -8270 1995
rect -8250 1975 -8180 1995
rect -8160 1975 -8135 1995
rect -8115 1975 -8090 1995
rect -8070 1975 -8000 1995
rect -7980 1975 -7955 1995
rect -7935 1975 -7910 1995
rect -7890 1975 -7820 1995
rect -7800 1975 -7775 1995
rect -7755 1975 -7730 1995
rect -7710 1975 -7640 1995
rect -7620 1975 -7595 1995
rect -7575 1975 -7550 1995
rect -7530 1975 -7460 1995
rect -7440 1975 -7415 1995
rect -7395 1975 -7370 1995
rect -7350 1975 -7280 1995
rect -7260 1975 -7235 1995
rect -7215 1975 -7190 1995
rect -7170 1975 -7100 1995
rect -7080 1975 -7055 1995
rect -7035 1975 -7010 1995
rect -6990 1975 -6920 1995
rect -6900 1975 -6875 1995
rect -6855 1975 -6830 1995
rect -6810 1975 -6740 1995
rect -6720 1975 -6695 1995
rect -6675 1975 -6650 1995
rect -6630 1975 -6560 1995
rect -6540 1975 -6515 1995
rect -6495 1975 -6470 1995
rect -6450 1975 -6380 1995
rect -6360 1975 -6335 1995
rect -6315 1975 -6290 1995
rect -6270 1975 -6200 1995
rect -6180 1975 -6155 1995
rect -6135 1975 -6110 1995
rect -6090 1975 -6020 1995
rect -6000 1975 -5975 1995
rect -5955 1975 -5930 1995
rect -5910 1975 -5840 1995
rect -5820 1975 -5795 1995
rect -5775 1975 -5750 1995
rect -5730 1975 -5660 1995
rect -5640 1975 -5615 1995
rect -5595 1975 -5570 1995
rect -5550 1975 -5480 1995
rect -5460 1975 -5435 1995
rect -5415 1975 -5390 1995
rect -5370 1975 -5300 1995
rect -5280 1975 -5255 1995
rect -5235 1975 -5210 1995
rect -5190 1975 -5120 1995
rect -5100 1975 -5075 1995
rect -5055 1975 -5030 1995
rect -5010 1975 -4940 1995
rect -4920 1975 -4895 1995
rect -4875 1975 -4850 1995
rect -4830 1975 -4760 1995
rect -4740 1975 -4715 1995
rect -4695 1975 -4670 1995
rect -4650 1975 -4580 1995
rect -4560 1975 -4535 1995
rect -4515 1975 -4490 1995
rect -4470 1975 -4400 1995
rect -4380 1975 -4355 1995
rect -4335 1975 -4310 1995
rect -4290 1975 -4220 1995
rect -4200 1975 -4175 1995
rect -4155 1975 -4130 1995
rect -4110 1975 -4040 1995
rect -4020 1975 -3995 1995
rect -3975 1975 -3950 1995
rect -3930 1975 -3860 1995
rect -3840 1975 -3815 1995
rect -3795 1975 -3770 1995
rect -3750 1975 -3680 1995
rect -3660 1975 -3635 1995
rect -3615 1975 -3590 1995
rect -3570 1975 -3500 1995
rect -3480 1975 -3455 1995
rect -3435 1975 -3410 1995
rect -3390 1975 -3320 1995
rect -3300 1975 -3275 1995
rect -3255 1975 -3230 1995
rect -3210 1975 -3140 1995
rect -3120 1975 -3095 1995
rect -3075 1975 -3050 1995
rect -3030 1975 -2960 1995
rect -2940 1975 -2915 1995
rect -2895 1975 -2870 1995
rect -2850 1975 -2780 1995
rect -2760 1975 -2735 1995
rect -2715 1975 -2690 1995
rect -2670 1975 -2600 1995
rect -2580 1975 -2555 1995
rect -2535 1975 -2510 1995
rect -2490 1975 -2420 1995
rect -2400 1975 -2375 1995
rect -2355 1975 -2330 1995
rect -2310 1975 -2240 1995
rect -2220 1975 -2195 1995
rect -2175 1975 -2150 1995
rect -2130 1975 -2060 1995
rect -2040 1975 -2015 1995
rect -1995 1975 -1970 1995
rect -1950 1975 -1880 1995
rect -1860 1975 -1835 1995
rect -1815 1975 -1790 1995
rect -1770 1975 -1700 1995
rect -1680 1975 -1655 1995
rect -1635 1975 -1610 1995
rect -1590 1975 -1520 1995
rect -1500 1975 -1475 1995
rect -1455 1975 -1430 1995
rect -1410 1975 -1340 1995
rect -1320 1975 -1295 1995
rect -1275 1975 -1250 1995
rect -1230 1975 -1160 1995
rect -1140 1975 -1115 1995
rect -1095 1975 -1070 1995
rect -1050 1975 -980 1995
rect -960 1975 -935 1995
rect -915 1975 -890 1995
rect -870 1975 -800 1995
rect -780 1975 -755 1995
rect -735 1975 -710 1995
rect -690 1975 -620 1995
rect -600 1975 -530 1995
rect -510 1975 -440 1995
rect -420 1975 -350 1995
rect -330 1975 -260 1995
rect -240 1975 -170 1995
rect -150 1975 -80 1995
rect -60 1975 -35 1995
rect -15 1975 100 1995
rect 120 1975 130 1995
rect -11690 1775 -11670 1975
rect -11555 1935 -11535 1945
rect -11555 1845 -11535 1855
rect -11465 1935 -11445 1945
rect -11465 1845 -11445 1855
rect -11375 1935 -11355 1945
rect -11375 1845 -11355 1855
rect -11285 1935 -11265 1945
rect -11285 1820 -11265 1855
rect -11195 1935 -11175 1945
rect -11195 1845 -11175 1855
rect -11105 1935 -11085 1945
rect -11105 1820 -11085 1855
rect -11015 1935 -10995 1945
rect -11015 1845 -10995 1855
rect -10925 1935 -10905 1945
rect -10925 1845 -10905 1855
rect -10835 1935 -10815 1945
rect -10835 1845 -10815 1855
rect -10745 1935 -10725 1945
rect -10745 1845 -10725 1855
rect -10655 1935 -10635 1945
rect -10655 1845 -10635 1855
rect -10565 1935 -10545 1945
rect -10565 1845 -10545 1855
rect -10475 1935 -10455 1945
rect -10475 1845 -10455 1855
rect -10385 1935 -10365 1945
rect -10385 1845 -10365 1855
rect -10295 1935 -10275 1945
rect -10295 1845 -10275 1855
rect -10205 1935 -10185 1945
rect -10205 1845 -10185 1855
rect -10115 1935 -10095 1945
rect -10115 1845 -10095 1855
rect -10025 1935 -10005 1945
rect -10025 1845 -10005 1855
rect -9935 1935 -9915 1945
rect -9935 1845 -9915 1855
rect -9845 1935 -9825 1945
rect -9845 1845 -9825 1855
rect -9755 1935 -9735 1945
rect -9755 1845 -9735 1855
rect -9665 1935 -9645 1945
rect -9665 1845 -9645 1855
rect -9575 1935 -9555 1945
rect -9575 1845 -9555 1855
rect -9485 1935 -9465 1945
rect -9485 1845 -9465 1855
rect -9395 1935 -9375 1945
rect -9395 1845 -9375 1855
rect -9305 1935 -9285 1945
rect -9305 1845 -9285 1855
rect -9215 1935 -9195 1945
rect -9215 1845 -9195 1855
rect -9125 1935 -9105 1945
rect -9125 1845 -9105 1855
rect -9035 1935 -9015 1945
rect -9035 1845 -9015 1855
rect -8945 1935 -8925 1945
rect -8945 1845 -8925 1855
rect -8855 1935 -8835 1945
rect -8855 1845 -8835 1855
rect -8765 1935 -8745 1945
rect -8765 1845 -8745 1855
rect -8675 1935 -8655 1945
rect -8675 1845 -8655 1855
rect -8585 1935 -8565 1945
rect -8585 1845 -8565 1855
rect -8495 1935 -8475 1945
rect -8495 1845 -8475 1855
rect -8405 1935 -8385 1945
rect -8405 1845 -8385 1855
rect -8315 1935 -8295 1945
rect -8315 1845 -8295 1855
rect -8225 1935 -8205 1945
rect -8225 1845 -8205 1855
rect -8135 1935 -8115 1945
rect -8135 1845 -8115 1855
rect -8045 1935 -8025 1945
rect -8045 1845 -8025 1855
rect -7955 1935 -7935 1945
rect -7955 1845 -7935 1855
rect -7865 1935 -7845 1945
rect -7865 1845 -7845 1855
rect -7775 1935 -7755 1945
rect -7775 1845 -7755 1855
rect -7685 1935 -7665 1945
rect -7685 1845 -7665 1855
rect -7595 1935 -7575 1945
rect -7595 1845 -7575 1855
rect -7505 1935 -7485 1945
rect -7505 1845 -7485 1855
rect -7415 1935 -7395 1945
rect -7415 1845 -7395 1855
rect -7325 1935 -7305 1945
rect -7325 1845 -7305 1855
rect -7235 1935 -7215 1945
rect -7235 1845 -7215 1855
rect -7145 1935 -7125 1945
rect -7145 1845 -7125 1855
rect -7055 1935 -7035 1945
rect -7055 1845 -7035 1855
rect -6965 1935 -6945 1945
rect -6965 1845 -6945 1855
rect -6875 1935 -6855 1945
rect -6875 1845 -6855 1855
rect -6785 1935 -6765 1945
rect -6785 1845 -6765 1855
rect -6695 1935 -6675 1945
rect -6695 1845 -6675 1855
rect -6605 1935 -6585 1945
rect -6605 1845 -6585 1855
rect -6515 1935 -6495 1945
rect -6515 1845 -6495 1855
rect -6425 1935 -6405 1945
rect -6425 1845 -6405 1855
rect -6335 1935 -6315 1945
rect -6335 1845 -6315 1855
rect -6245 1935 -6225 1945
rect -6245 1845 -6225 1855
rect -6155 1935 -6135 1945
rect -6155 1820 -6135 1855
rect -6065 1935 -6045 1945
rect -6065 1845 -6045 1855
rect -5975 1935 -5955 1945
rect -5975 1845 -5955 1855
rect -5885 1935 -5865 1945
rect -5885 1845 -5865 1855
rect -5795 1935 -5775 1945
rect -5795 1845 -5775 1855
rect -5705 1935 -5685 1945
rect -5705 1845 -5685 1855
rect -5615 1935 -5595 1945
rect -5615 1845 -5595 1855
rect -5525 1935 -5505 1945
rect -5525 1845 -5505 1855
rect -5435 1935 -5415 1945
rect -5435 1845 -5415 1855
rect -5345 1935 -5325 1945
rect -5345 1845 -5325 1855
rect -5255 1935 -5235 1945
rect -5255 1845 -5235 1855
rect -5165 1935 -5145 1945
rect -5165 1845 -5145 1855
rect -5075 1935 -5055 1945
rect -5075 1845 -5055 1855
rect -4985 1935 -4965 1945
rect -4985 1845 -4965 1855
rect -4895 1935 -4875 1945
rect -4895 1845 -4875 1855
rect -4805 1935 -4785 1945
rect -4805 1845 -4785 1855
rect -4715 1935 -4695 1945
rect -4715 1845 -4695 1855
rect -4625 1935 -4605 1945
rect -4625 1845 -4605 1855
rect -4535 1935 -4515 1945
rect -4535 1845 -4515 1855
rect -4445 1935 -4425 1945
rect -4445 1845 -4425 1855
rect -4355 1935 -4335 1945
rect -4355 1845 -4335 1855
rect -4265 1935 -4245 1945
rect -4265 1845 -4245 1855
rect -4175 1935 -4155 1945
rect -4175 1845 -4155 1855
rect -4085 1935 -4065 1945
rect -4085 1845 -4065 1855
rect -3995 1935 -3975 1945
rect -3995 1845 -3975 1855
rect -3905 1935 -3885 1945
rect -3905 1845 -3885 1855
rect -3815 1935 -3795 1945
rect -3815 1845 -3795 1855
rect -3725 1935 -3705 1945
rect -3725 1845 -3705 1855
rect -3635 1935 -3615 1945
rect -3635 1845 -3615 1855
rect -3545 1935 -3525 1945
rect -3545 1845 -3525 1855
rect -3455 1935 -3435 1945
rect -3455 1845 -3435 1855
rect -3365 1935 -3345 1945
rect -3365 1845 -3345 1855
rect -3275 1935 -3255 1945
rect -3275 1845 -3255 1855
rect -3185 1935 -3165 1945
rect -3185 1845 -3165 1855
rect -3095 1935 -3075 1945
rect -3095 1845 -3075 1855
rect -3005 1935 -2985 1945
rect -3005 1845 -2985 1855
rect -2915 1935 -2895 1945
rect -2915 1845 -2895 1855
rect -2825 1935 -2805 1945
rect -2825 1845 -2805 1855
rect -2735 1935 -2715 1945
rect -2735 1845 -2715 1855
rect -2645 1935 -2625 1945
rect -2645 1845 -2625 1855
rect -2555 1935 -2535 1945
rect -2555 1820 -2535 1855
rect -2465 1935 -2445 1945
rect -2465 1845 -2445 1855
rect -2375 1935 -2355 1945
rect -2375 1845 -2355 1855
rect -2285 1935 -2265 1945
rect -2285 1845 -2265 1855
rect -2195 1935 -2175 1945
rect -2195 1845 -2175 1855
rect -2105 1935 -2085 1945
rect -2105 1845 -2085 1855
rect -2015 1935 -1995 1945
rect -2015 1845 -1995 1855
rect -1925 1935 -1905 1945
rect -1925 1845 -1905 1855
rect -1835 1935 -1815 1945
rect -1835 1845 -1815 1855
rect -1745 1935 -1725 1945
rect -1745 1845 -1725 1855
rect -1655 1935 -1635 1945
rect -1655 1845 -1635 1855
rect -1565 1935 -1545 1945
rect -1565 1845 -1545 1855
rect -1475 1935 -1455 1945
rect -1475 1845 -1455 1855
rect -1385 1935 -1365 1945
rect -1385 1845 -1365 1855
rect -1295 1935 -1275 1945
rect -1295 1845 -1275 1855
rect -1205 1935 -1185 1945
rect -1205 1845 -1185 1855
rect -1115 1935 -1095 1945
rect -1115 1845 -1095 1855
rect -1025 1935 -1005 1945
rect -1025 1845 -1005 1855
rect -935 1935 -915 1945
rect -935 1845 -915 1855
rect -845 1935 -825 1945
rect -845 1845 -825 1855
rect -755 1935 -735 1945
rect -755 1845 -735 1855
rect -665 1935 -645 1945
rect -665 1845 -645 1855
rect -575 1935 -555 1945
rect -575 1845 -555 1855
rect -485 1935 -465 1945
rect -485 1820 -465 1855
rect -395 1935 -375 1945
rect -395 1845 -375 1855
rect -305 1935 -285 1945
rect -305 1820 -285 1855
rect -215 1935 -195 1945
rect -215 1845 -195 1855
rect -125 1935 -105 1945
rect -125 1845 -105 1855
rect -35 1935 -15 1945
rect -35 1845 -15 1855
rect -11520 1800 -11510 1820
rect -11490 1800 -11420 1820
rect -11400 1800 -11330 1820
rect -11310 1800 -11240 1820
rect -11220 1800 -11150 1820
rect -11130 1800 -11060 1820
rect -11040 1800 -10970 1820
rect -10950 1800 -10880 1820
rect -10860 1800 -10850 1820
rect -10800 1800 -10790 1820
rect -10770 1800 -10700 1820
rect -10680 1800 -10670 1820
rect -10620 1800 -10610 1820
rect -10590 1800 -10520 1820
rect -10500 1800 -10490 1820
rect -10440 1800 -10430 1820
rect -10410 1800 -10340 1820
rect -10320 1800 -10310 1820
rect -10260 1800 -10250 1820
rect -10230 1800 -10160 1820
rect -10140 1800 -10130 1820
rect -10080 1800 -10070 1820
rect -10050 1800 -9980 1820
rect -9960 1800 -9950 1820
rect -9900 1800 -9890 1820
rect -9870 1800 -9800 1820
rect -9780 1800 -9770 1820
rect -9720 1800 -9710 1820
rect -9690 1800 -9620 1820
rect -9600 1800 -9590 1820
rect -9540 1800 -9530 1820
rect -9510 1800 -9440 1820
rect -9420 1800 -9410 1820
rect -9360 1800 -9350 1820
rect -9330 1800 -9260 1820
rect -9240 1800 -9230 1820
rect -9180 1800 -9170 1820
rect -9150 1800 -9080 1820
rect -9060 1800 -9050 1820
rect -9000 1800 -8990 1820
rect -8970 1800 -8900 1820
rect -8880 1800 -8870 1820
rect -8820 1800 -8810 1820
rect -8790 1800 -8720 1820
rect -8700 1800 -8690 1820
rect -8640 1800 -8630 1820
rect -8610 1800 -8540 1820
rect -8520 1800 -8510 1820
rect -8460 1800 -8450 1820
rect -8430 1800 -8360 1820
rect -8340 1800 -8330 1820
rect -8280 1800 -8270 1820
rect -8250 1800 -8180 1820
rect -8160 1800 -8150 1820
rect -8100 1800 -8090 1820
rect -8070 1800 -8000 1820
rect -7980 1800 -7970 1820
rect -7920 1800 -7910 1820
rect -7890 1800 -7820 1820
rect -7800 1800 -7790 1820
rect -7740 1800 -7730 1820
rect -7710 1800 -7640 1820
rect -7620 1800 -7610 1820
rect -7560 1800 -7550 1820
rect -7530 1800 -7460 1820
rect -7440 1800 -7430 1820
rect -7380 1800 -7370 1820
rect -7350 1800 -7280 1820
rect -7260 1800 -7250 1820
rect -7200 1800 -7190 1820
rect -7170 1800 -7100 1820
rect -7080 1800 -7010 1820
rect -6990 1800 -6920 1820
rect -6900 1800 -6830 1820
rect -6810 1800 -6740 1820
rect -6720 1800 -6650 1820
rect -6630 1800 -6560 1820
rect -6540 1800 -6470 1820
rect -6450 1800 -6380 1820
rect -6360 1800 -6290 1820
rect -6270 1800 -6200 1820
rect -6180 1800 -6110 1820
rect -6090 1800 -6020 1820
rect -6000 1800 -5930 1820
rect -5910 1800 -5840 1820
rect -5820 1800 -5750 1820
rect -5730 1800 -5660 1820
rect -5640 1800 -5570 1820
rect -5550 1800 -5480 1820
rect -5460 1800 -5390 1820
rect -5370 1800 -5300 1820
rect -5280 1800 -5210 1820
rect -5190 1800 -5120 1820
rect -5100 1800 -5090 1820
rect -5040 1800 -5030 1820
rect -5010 1800 -4940 1820
rect -4920 1800 -4910 1820
rect -4860 1800 -4850 1820
rect -4830 1800 -4760 1820
rect -4740 1800 -4730 1820
rect -4680 1800 -4670 1820
rect -4650 1800 -4580 1820
rect -4560 1800 -4550 1820
rect -4500 1800 -4490 1820
rect -4470 1800 -4400 1820
rect -4380 1800 -4370 1820
rect -4320 1800 -4310 1820
rect -4290 1800 -4220 1820
rect -4200 1800 -4190 1820
rect -4140 1800 -4130 1820
rect -4110 1800 -4040 1820
rect -4020 1800 -4010 1820
rect -3960 1800 -3950 1820
rect -3930 1800 -3860 1820
rect -3840 1800 -3830 1820
rect -3780 1800 -3770 1820
rect -3750 1800 -3680 1820
rect -3660 1800 -3650 1820
rect -3600 1800 -3590 1820
rect -3570 1800 -3500 1820
rect -3480 1800 -3410 1820
rect -3390 1800 -3320 1820
rect -3300 1800 -3230 1820
rect -3210 1800 -3140 1820
rect -3120 1800 -3050 1820
rect -3030 1800 -2960 1820
rect -2940 1800 -2870 1820
rect -2850 1800 -2780 1820
rect -2760 1800 -2690 1820
rect -2670 1800 -2600 1820
rect -2580 1800 -2510 1820
rect -2490 1800 -2420 1820
rect -2400 1800 -2330 1820
rect -2310 1800 -2240 1820
rect -2220 1800 -2150 1820
rect -2130 1800 -2060 1820
rect -2040 1800 -1970 1820
rect -1950 1800 -1880 1820
rect -1860 1800 -1790 1820
rect -1770 1800 -1700 1820
rect -1680 1800 -1610 1820
rect -1590 1800 -1520 1820
rect -1500 1800 -1490 1820
rect -1440 1800 -1430 1820
rect -1410 1800 -1340 1820
rect -1320 1800 -1310 1820
rect -1260 1800 -1250 1820
rect -1230 1800 -1160 1820
rect -1140 1800 -1130 1820
rect -1080 1800 -1070 1820
rect -1050 1800 -980 1820
rect -960 1800 -950 1820
rect -900 1800 -890 1820
rect -870 1800 -800 1820
rect -780 1800 -770 1820
rect -720 1800 -710 1820
rect -690 1800 -620 1820
rect -600 1800 -530 1820
rect -510 1800 -440 1820
rect -420 1800 -350 1820
rect -330 1800 -260 1820
rect -240 1800 -170 1820
rect -150 1800 -80 1820
rect -60 1800 -50 1820
rect 100 1775 120 1975
rect -11690 1755 -11510 1775
rect -11490 1755 -11420 1775
rect -11400 1755 -11330 1775
rect -11310 1755 -11240 1775
rect -11220 1755 -11150 1775
rect -11130 1755 -11060 1775
rect -11040 1755 -10970 1775
rect -10950 1755 -10880 1775
rect -10860 1755 -10790 1775
rect -10770 1755 -10700 1775
rect -10680 1755 -10610 1775
rect -10590 1755 -10520 1775
rect -10500 1755 -10430 1775
rect -10410 1755 -10340 1775
rect -10320 1755 -10250 1775
rect -10230 1755 -10160 1775
rect -10140 1755 -10070 1775
rect -10050 1755 -9980 1775
rect -9960 1755 -9890 1775
rect -9870 1755 -9800 1775
rect -9780 1755 -9710 1775
rect -9690 1755 -9620 1775
rect -9600 1755 -9530 1775
rect -9510 1755 -9440 1775
rect -9420 1755 -9350 1775
rect -9330 1755 -9260 1775
rect -9240 1755 -9170 1775
rect -9150 1755 -9080 1775
rect -9060 1755 -8990 1775
rect -8970 1755 -8900 1775
rect -8880 1755 -8810 1775
rect -8790 1755 -8720 1775
rect -8700 1755 -8630 1775
rect -8610 1755 -8540 1775
rect -8520 1755 -8450 1775
rect -8430 1755 -8360 1775
rect -8340 1755 -8270 1775
rect -8250 1755 -8180 1775
rect -8160 1755 -8090 1775
rect -8070 1755 -8000 1775
rect -7980 1755 -7910 1775
rect -7890 1755 -7820 1775
rect -7800 1755 -7730 1775
rect -7710 1755 -7640 1775
rect -7620 1755 -7550 1775
rect -7530 1755 -7460 1775
rect -7440 1755 -7370 1775
rect -7350 1755 -7280 1775
rect -7260 1755 -7190 1775
rect -7170 1755 -7100 1775
rect -7080 1755 -7010 1775
rect -6990 1755 -6920 1775
rect -6900 1755 -6830 1775
rect -6810 1755 -6740 1775
rect -6720 1755 -6650 1775
rect -6630 1755 -6560 1775
rect -6540 1755 -6470 1775
rect -6450 1755 -6380 1775
rect -6360 1755 -6290 1775
rect -6270 1755 -6200 1775
rect -6180 1755 -6110 1775
rect -6090 1755 -6020 1775
rect -6000 1755 -5930 1775
rect -5910 1755 -5840 1775
rect -5820 1755 -5750 1775
rect -5730 1755 -5660 1775
rect -5640 1755 -5570 1775
rect -5550 1755 -5480 1775
rect -5460 1755 -5390 1775
rect -5370 1755 -5300 1775
rect -5280 1755 -5210 1775
rect -5190 1755 -5120 1775
rect -5100 1755 -5030 1775
rect -5010 1755 -4940 1775
rect -4920 1755 -4850 1775
rect -4830 1755 -4760 1775
rect -4740 1755 -4670 1775
rect -4650 1755 -4580 1775
rect -4560 1755 -4490 1775
rect -4470 1755 -4400 1775
rect -4380 1755 -4310 1775
rect -4290 1755 -4220 1775
rect -4200 1755 -4130 1775
rect -4110 1755 -4040 1775
rect -4020 1755 -3950 1775
rect -3930 1755 -3860 1775
rect -3840 1755 -3770 1775
rect -3750 1755 -3680 1775
rect -3660 1755 -3590 1775
rect -3570 1755 -3500 1775
rect -3480 1755 -3410 1775
rect -3390 1755 -3320 1775
rect -3300 1755 -3230 1775
rect -3210 1755 -3140 1775
rect -3120 1755 -3050 1775
rect -3030 1755 -2960 1775
rect -2940 1755 -2870 1775
rect -2850 1755 -2780 1775
rect -2760 1755 -2690 1775
rect -2670 1755 -2600 1775
rect -2580 1755 -2510 1775
rect -2490 1755 -2420 1775
rect -2400 1755 -2330 1775
rect -2310 1755 -2240 1775
rect -2220 1755 -2150 1775
rect -2130 1755 -2060 1775
rect -2040 1755 -1970 1775
rect -1950 1755 -1880 1775
rect -1860 1755 -1790 1775
rect -1770 1755 -1700 1775
rect -1680 1755 -1610 1775
rect -1590 1755 -1520 1775
rect -1500 1755 -1430 1775
rect -1410 1755 -1340 1775
rect -1320 1755 -1250 1775
rect -1230 1755 -1160 1775
rect -1140 1755 -1070 1775
rect -1050 1755 -980 1775
rect -960 1755 -890 1775
rect -870 1755 -800 1775
rect -780 1755 -710 1775
rect -690 1755 -620 1775
rect -600 1755 -530 1775
rect -510 1755 -440 1775
rect -420 1755 -350 1775
rect -330 1755 -260 1775
rect -240 1755 -170 1775
rect -150 1755 -80 1775
rect -60 1755 120 1775
rect -11565 1715 -10700 1735
rect -10680 1715 -10520 1735
rect -10500 1715 -9620 1735
rect -9600 1715 -9440 1735
rect -9420 1715 -9260 1735
rect -9240 1715 -9080 1735
rect -9060 1715 -8180 1735
rect -8160 1715 -8000 1735
rect -7980 1715 -7820 1735
rect -7800 1715 -7640 1735
rect -7620 1715 -4580 1735
rect -4560 1715 -4400 1735
rect -4380 1715 -4220 1735
rect -4200 1715 -4040 1735
rect -4020 1715 -980 1735
rect -960 1715 -800 1735
rect -780 1715 -125 1735
rect -105 1715 -5 1735
rect -11565 1675 -10340 1695
rect -10320 1675 -10160 1695
rect -10140 1675 -9980 1695
rect -9960 1675 -9800 1695
rect -9780 1675 -8900 1695
rect -8880 1675 -8720 1695
rect -8700 1675 -8540 1695
rect -8520 1675 -8360 1695
rect -8340 1675 -7460 1695
rect -7440 1675 -7280 1695
rect -7260 1675 -4940 1695
rect -4920 1675 -4760 1695
rect -4740 1675 -3860 1695
rect -3840 1675 -3680 1695
rect -3660 1675 -1340 1695
rect -1320 1675 -1160 1695
rect -1140 1675 -215 1695
rect -195 1675 -5 1695
rect -11565 1635 -11105 1655
rect -11085 1635 -9035 1655
rect -9015 1635 -8315 1655
rect -8295 1635 -3995 1655
rect -3975 1635 -3545 1655
rect -3525 1635 -3365 1655
rect -3345 1635 -3185 1655
rect -3165 1635 -3005 1655
rect -2985 1635 -2825 1655
rect -2805 1635 -2645 1655
rect -2625 1635 -2465 1655
rect -2445 1635 -2285 1655
rect -2265 1635 -2105 1655
rect -2085 1635 -1925 1655
rect -1905 1635 -1745 1655
rect -1725 1635 -1565 1655
rect -1545 1635 -1115 1655
rect -1095 1635 -5 1655
rect -11565 1595 -11195 1615
rect -11175 1595 -10475 1615
rect -10455 1595 -9755 1615
rect -9735 1595 -7595 1615
rect -7575 1595 -7145 1615
rect -7125 1595 -6965 1615
rect -6945 1595 -6785 1615
rect -6765 1595 -6605 1615
rect -6585 1595 -6425 1615
rect -6405 1595 -6245 1615
rect -6225 1595 -6065 1615
rect -6045 1595 -5885 1615
rect -5865 1595 -5705 1615
rect -5685 1595 -5525 1615
rect -5505 1595 -5345 1615
rect -5325 1595 -5165 1615
rect -5145 1595 -4715 1615
rect -4695 1595 -5 1615
rect -11565 1555 -11285 1575
rect -11265 1555 -3590 1575
rect -3570 1555 -3410 1575
rect -3390 1555 -3230 1575
rect -3210 1555 -3050 1575
rect -3030 1555 -2870 1575
rect -2850 1555 -2690 1575
rect -2670 1555 -2510 1575
rect -2490 1555 -2330 1575
rect -2310 1555 -2150 1575
rect -2130 1555 -1970 1575
rect -1950 1555 -1790 1575
rect -1770 1555 -1610 1575
rect -1590 1555 -5 1575
rect -11565 1515 -11375 1535
rect -11355 1515 -7190 1535
rect -7170 1515 -7010 1535
rect -6990 1515 -6830 1535
rect -6810 1515 -6650 1535
rect -6630 1515 -6470 1535
rect -6450 1515 -6290 1535
rect -6270 1515 -6110 1535
rect -6090 1515 -5930 1535
rect -5910 1515 -5750 1535
rect -5730 1515 -5570 1535
rect -5550 1515 -5390 1535
rect -5370 1515 -5210 1535
rect -5190 1515 -5 1535
rect -11565 1475 -11465 1495
rect -11445 1475 -10115 1495
rect -10095 1475 -7235 1495
rect -7215 1475 -5075 1495
rect -5055 1475 -5 1495
rect -11565 1435 -10790 1455
rect -10770 1435 -10610 1455
rect -10590 1435 -9710 1455
rect -9690 1435 -9530 1455
rect -9510 1435 -9350 1455
rect -9330 1435 -9170 1455
rect -9150 1435 -8675 1455
rect -8655 1435 -8270 1455
rect -8250 1435 -8090 1455
rect -8070 1435 -3635 1455
rect -3615 1435 -1475 1455
rect -1455 1435 -485 1455
rect -465 1435 -5 1455
rect -11565 1395 -10430 1415
rect -10410 1395 -10250 1415
rect -10230 1395 -10070 1415
rect -10050 1395 -9890 1415
rect -9870 1395 -8990 1415
rect -8970 1395 -8810 1415
rect -8790 1395 -8630 1415
rect -8610 1395 -8450 1415
rect -8430 1395 -7550 1415
rect -7530 1395 -7370 1415
rect -7350 1395 -5030 1415
rect -5010 1395 -4850 1415
rect -4830 1395 -3950 1415
rect -3930 1395 -3770 1415
rect -3750 1395 -1430 1415
rect -1410 1395 -1250 1415
rect -1230 1395 -305 1415
rect -285 1395 -5 1415
rect -11565 1355 -7910 1375
rect -7890 1355 -7730 1375
rect -7710 1355 -4670 1375
rect -4650 1355 -4490 1375
rect -4470 1355 -4310 1375
rect -4290 1355 -4130 1375
rect -4110 1355 -1070 1375
rect -1050 1355 -890 1375
rect -870 1355 -395 1375
rect -375 1355 -5 1375
rect -11690 1315 -11510 1335
rect -11490 1315 -11420 1335
rect -11400 1315 -11330 1335
rect -11310 1315 -11240 1335
rect -11220 1315 -11150 1335
rect -11130 1315 -11060 1335
rect -11040 1315 -10970 1335
rect -10950 1315 -10880 1335
rect -10860 1315 -10790 1335
rect -10770 1315 -10700 1335
rect -10680 1315 -10610 1335
rect -10590 1315 -10520 1335
rect -10500 1315 -10430 1335
rect -10410 1315 -10340 1335
rect -10320 1315 -10250 1335
rect -10230 1315 -10160 1335
rect -10140 1315 -10070 1335
rect -10050 1315 -9980 1335
rect -9960 1315 -9890 1335
rect -9870 1315 -9800 1335
rect -9780 1315 -9710 1335
rect -9690 1315 -9620 1335
rect -9600 1315 -9530 1335
rect -9510 1315 -9440 1335
rect -9420 1315 -9350 1335
rect -9330 1315 -9260 1335
rect -9240 1315 -9170 1335
rect -9150 1315 -9080 1335
rect -9060 1315 -8990 1335
rect -8970 1315 -8900 1335
rect -8880 1315 -8810 1335
rect -8790 1315 -8720 1335
rect -8700 1315 -8630 1335
rect -8610 1315 -8540 1335
rect -8520 1315 -8450 1335
rect -8430 1315 -8360 1335
rect -8340 1315 -8270 1335
rect -8250 1315 -8180 1335
rect -8160 1315 -8090 1335
rect -8070 1315 -8000 1335
rect -7980 1315 -7910 1335
rect -7890 1315 -7820 1335
rect -7800 1315 -7730 1335
rect -7710 1315 -7640 1335
rect -7620 1315 -7550 1335
rect -7530 1315 -7460 1335
rect -7440 1315 -7370 1335
rect -7350 1315 -7280 1335
rect -7260 1315 -7190 1335
rect -7170 1315 -7100 1335
rect -7080 1315 -7010 1335
rect -6990 1315 -6920 1335
rect -6900 1315 -6830 1335
rect -6810 1315 -6740 1335
rect -6720 1315 -6650 1335
rect -6630 1315 -6560 1335
rect -6540 1315 -6470 1335
rect -6450 1315 -6380 1335
rect -6360 1315 -6290 1335
rect -6270 1315 -6200 1335
rect -6180 1315 -6110 1335
rect -6090 1315 -6020 1335
rect -6000 1315 -5930 1335
rect -5910 1315 -5840 1335
rect -5820 1315 -5750 1335
rect -5730 1315 -5660 1335
rect -5640 1315 -5570 1335
rect -5550 1315 -5480 1335
rect -5460 1315 -5390 1335
rect -5370 1315 -5300 1335
rect -5280 1315 -5210 1335
rect -5190 1315 -5120 1335
rect -5100 1315 -5030 1335
rect -5010 1315 -4940 1335
rect -4920 1315 -4850 1335
rect -4830 1315 -4760 1335
rect -4740 1315 -4670 1335
rect -4650 1315 -4580 1335
rect -4560 1315 -4490 1335
rect -4470 1315 -4400 1335
rect -4380 1315 -4310 1335
rect -4290 1315 -4220 1335
rect -4200 1315 -4130 1335
rect -4110 1315 -4040 1335
rect -4020 1315 -3950 1335
rect -3930 1315 -3860 1335
rect -3840 1315 -3770 1335
rect -3750 1315 -3680 1335
rect -3660 1315 -3590 1335
rect -3570 1315 -3500 1335
rect -3480 1315 -3410 1335
rect -3390 1315 -3320 1335
rect -3300 1315 -3230 1335
rect -3210 1315 -3140 1335
rect -3120 1315 -3050 1335
rect -3030 1315 -2960 1335
rect -2940 1315 -2870 1335
rect -2850 1315 -2780 1335
rect -2760 1315 -2690 1335
rect -2670 1315 -2600 1335
rect -2580 1315 -2510 1335
rect -2490 1315 -2420 1335
rect -2400 1315 -2330 1335
rect -2310 1315 -2240 1335
rect -2220 1315 -2150 1335
rect -2130 1315 -2060 1335
rect -2040 1315 -1970 1335
rect -1950 1315 -1880 1335
rect -1860 1315 -1790 1335
rect -1770 1315 -1700 1335
rect -1680 1315 -1610 1335
rect -1590 1315 -1520 1335
rect -1500 1315 -1430 1335
rect -1410 1315 -1340 1335
rect -1320 1315 -1250 1335
rect -1230 1315 -1160 1335
rect -1140 1315 -1070 1335
rect -1050 1315 -980 1335
rect -960 1315 -890 1335
rect -870 1315 -800 1335
rect -780 1315 -710 1335
rect -690 1315 -620 1335
rect -600 1315 -530 1335
rect -510 1315 -440 1335
rect -420 1315 -350 1335
rect -330 1315 -260 1335
rect -240 1315 -170 1335
rect -150 1315 -80 1335
rect -60 1315 120 1335
rect -11690 680 -11670 1315
rect -11565 1275 -7235 1295
rect -7215 1275 -7055 1295
rect -7035 1275 -6875 1295
rect -6855 1275 -6695 1295
rect -6675 1275 -6515 1295
rect -6495 1275 -6335 1295
rect -6315 1275 -6155 1295
rect -6135 1275 -5975 1295
rect -5955 1275 -5795 1295
rect -5775 1275 -5615 1295
rect -5595 1275 -5435 1295
rect -5415 1275 -5255 1295
rect -5235 1275 -5075 1295
rect -5055 1275 -3635 1295
rect -3615 1275 -3455 1295
rect -3435 1275 -3275 1295
rect -3255 1275 -3095 1295
rect -3075 1275 -2915 1295
rect -2895 1275 -2735 1295
rect -2715 1275 -2555 1295
rect -2535 1275 -2375 1295
rect -2355 1275 -2195 1295
rect -2175 1275 -2015 1295
rect -1995 1275 -1835 1295
rect -1815 1275 -1655 1295
rect -1635 1275 -1475 1295
rect -1455 1275 -575 1295
rect -555 1275 -5 1295
rect -11615 1235 -11510 1255
rect -11490 1235 -11420 1255
rect -11400 1235 -11330 1255
rect -11310 1235 -11240 1255
rect -11220 1235 -11150 1255
rect -11130 1235 -11060 1255
rect -11040 1235 -10970 1255
rect -10950 1235 -10880 1255
rect -10860 1235 -10790 1255
rect -10770 1235 -10700 1255
rect -10680 1235 -10610 1255
rect -10590 1235 -10520 1255
rect -10500 1235 -10430 1255
rect -10410 1235 -10340 1255
rect -10320 1235 -10250 1255
rect -10230 1235 -10160 1255
rect -10140 1235 -10070 1255
rect -10050 1235 -9980 1255
rect -9960 1235 -9890 1255
rect -9870 1235 -9800 1255
rect -9780 1235 -9710 1255
rect -9690 1235 -9620 1255
rect -9600 1235 -9530 1255
rect -9510 1235 -9440 1255
rect -9420 1235 -9350 1255
rect -9330 1235 -9260 1255
rect -9240 1235 -9170 1255
rect -9150 1235 -9080 1255
rect -9060 1235 -8990 1255
rect -8970 1235 -8900 1255
rect -8880 1235 -8810 1255
rect -8790 1235 -8720 1255
rect -8700 1235 -8630 1255
rect -8610 1235 -8540 1255
rect -8520 1235 -8450 1255
rect -8430 1235 -8360 1255
rect -8340 1235 -8270 1255
rect -8250 1235 -8180 1255
rect -8160 1235 -8090 1255
rect -8070 1235 -8000 1255
rect -7980 1235 -7910 1255
rect -7890 1235 -7820 1255
rect -7800 1235 -7730 1255
rect -7710 1235 -7640 1255
rect -7620 1235 -7550 1255
rect -7530 1235 -7460 1255
rect -7440 1235 -7370 1255
rect -7350 1235 -7280 1255
rect -7260 1235 -7190 1255
rect -7170 1235 -7100 1255
rect -7080 1235 -7010 1255
rect -6990 1235 -6920 1255
rect -6900 1235 -6830 1255
rect -6810 1235 -6740 1255
rect -6720 1235 -6650 1255
rect -6630 1235 -6560 1255
rect -6540 1235 -6470 1255
rect -6450 1235 -6380 1255
rect -6360 1235 -6290 1255
rect -6270 1235 -6200 1255
rect -6180 1235 -6110 1255
rect -6090 1235 -6020 1255
rect -6000 1235 -5930 1255
rect -5910 1235 -5840 1255
rect -5820 1235 -5750 1255
rect -5730 1235 -5660 1255
rect -5640 1235 -5570 1255
rect -5550 1235 -5480 1255
rect -5460 1235 -5390 1255
rect -5370 1235 -5300 1255
rect -5280 1235 -5210 1255
rect -5190 1235 -5120 1255
rect -5100 1235 -5030 1255
rect -5010 1235 -4940 1255
rect -4920 1235 -4850 1255
rect -4830 1235 -4760 1255
rect -4740 1235 -4670 1255
rect -4650 1235 -4580 1255
rect -4560 1235 -4490 1255
rect -4470 1235 -4400 1255
rect -4380 1235 -4310 1255
rect -4290 1235 -4220 1255
rect -4200 1235 -4130 1255
rect -4110 1235 -4040 1255
rect -4020 1235 -3950 1255
rect -3930 1235 -3860 1255
rect -3840 1235 -3770 1255
rect -3750 1235 -3680 1255
rect -3660 1235 -3590 1255
rect -3570 1235 -3500 1255
rect -3480 1235 -3410 1255
rect -3390 1235 -3320 1255
rect -3300 1235 -3230 1255
rect -3210 1235 -3140 1255
rect -3120 1235 -3050 1255
rect -3030 1235 -2960 1255
rect -2940 1235 -2870 1255
rect -2850 1235 -2780 1255
rect -2760 1235 -2690 1255
rect -2670 1235 -2600 1255
rect -2580 1235 -2510 1255
rect -2490 1235 -2420 1255
rect -2400 1235 -2330 1255
rect -2310 1235 -2240 1255
rect -2220 1235 -2150 1255
rect -2130 1235 -2060 1255
rect -2040 1235 -1970 1255
rect -1950 1235 -1880 1255
rect -1860 1235 -1790 1255
rect -1770 1235 -1700 1255
rect -1680 1235 -1610 1255
rect -1590 1235 -1520 1255
rect -1500 1235 -1430 1255
rect -1410 1235 -1340 1255
rect -1320 1235 -1250 1255
rect -1230 1235 -1160 1255
rect -1140 1235 -1070 1255
rect -1050 1235 -980 1255
rect -960 1235 -890 1255
rect -870 1235 -800 1255
rect -780 1235 -710 1255
rect -690 1235 -620 1255
rect -600 1235 -530 1255
rect -510 1235 -440 1255
rect -420 1235 -350 1255
rect -330 1235 -260 1255
rect -240 1235 -170 1255
rect -150 1235 -80 1255
rect -60 1235 45 1255
rect -11615 1035 -11595 1235
rect -11520 1190 -11510 1210
rect -11490 1190 -11420 1210
rect -11400 1190 -11330 1210
rect -11310 1190 -11240 1210
rect -11220 1190 -11150 1210
rect -11130 1190 -11060 1210
rect -11040 1190 -10970 1210
rect -10950 1190 -10880 1210
rect -10860 1190 -10845 1210
rect -10800 1190 -10790 1210
rect -10770 1190 -10700 1210
rect -10680 1190 -10670 1210
rect -10620 1190 -10610 1210
rect -10590 1190 -10520 1210
rect -10500 1190 -10490 1210
rect -10440 1190 -10430 1210
rect -10410 1190 -10340 1210
rect -10320 1190 -10310 1210
rect -10260 1190 -10250 1210
rect -10230 1190 -10160 1210
rect -10140 1190 -10130 1210
rect -10080 1190 -10070 1210
rect -10050 1190 -9980 1210
rect -9960 1190 -9950 1210
rect -9900 1190 -9890 1210
rect -9870 1190 -9800 1210
rect -9780 1190 -9770 1210
rect -9720 1190 -9710 1210
rect -9690 1190 -9620 1210
rect -9600 1190 -9590 1210
rect -9540 1190 -9530 1210
rect -9510 1190 -9440 1210
rect -9420 1190 -9410 1210
rect -9360 1190 -9350 1210
rect -9330 1190 -9260 1210
rect -9240 1190 -9230 1210
rect -9180 1190 -9170 1210
rect -9150 1190 -9080 1210
rect -9060 1190 -9050 1210
rect -9000 1190 -8990 1210
rect -8970 1190 -8900 1210
rect -8880 1190 -8870 1210
rect -8820 1190 -8810 1210
rect -8790 1190 -8720 1210
rect -8700 1190 -8690 1210
rect -8640 1190 -8630 1210
rect -8610 1190 -8540 1210
rect -8520 1190 -8510 1210
rect -8460 1190 -8450 1210
rect -8430 1190 -8360 1210
rect -8340 1190 -8330 1210
rect -8280 1190 -8270 1210
rect -8250 1190 -8180 1210
rect -8160 1190 -8150 1210
rect -8100 1190 -8090 1210
rect -8070 1190 -8000 1210
rect -7980 1190 -7970 1210
rect -7920 1190 -7910 1210
rect -7890 1190 -7820 1210
rect -7800 1190 -7790 1210
rect -7740 1190 -7730 1210
rect -7710 1190 -7640 1210
rect -7620 1190 -7610 1210
rect -7560 1190 -7550 1210
rect -7530 1190 -7460 1210
rect -7440 1190 -7430 1210
rect -7380 1190 -7370 1210
rect -7350 1190 -7280 1210
rect -7260 1190 -7250 1210
rect -7200 1190 -7190 1210
rect -7170 1190 -7100 1210
rect -7080 1190 -7070 1210
rect -7020 1190 -7010 1210
rect -6990 1190 -6920 1210
rect -6900 1190 -6890 1210
rect -6840 1190 -6830 1210
rect -6810 1190 -6740 1210
rect -6720 1190 -6710 1210
rect -6660 1190 -6650 1210
rect -6630 1190 -6560 1210
rect -6540 1190 -6530 1210
rect -6480 1190 -6470 1210
rect -6450 1190 -6380 1210
rect -6360 1190 -6350 1210
rect -6300 1190 -6290 1210
rect -6270 1190 -6200 1210
rect -6180 1190 -6170 1210
rect -6120 1190 -6110 1210
rect -6090 1190 -6020 1210
rect -6000 1190 -5990 1210
rect -5940 1190 -5930 1210
rect -5910 1190 -5840 1210
rect -5820 1190 -5810 1210
rect -5760 1190 -5750 1210
rect -5730 1190 -5660 1210
rect -5640 1190 -5630 1210
rect -5580 1190 -5570 1210
rect -5550 1190 -5480 1210
rect -5460 1190 -5450 1210
rect -5400 1190 -5390 1210
rect -5370 1190 -5300 1210
rect -5280 1190 -5270 1210
rect -5220 1190 -5210 1210
rect -5190 1190 -5120 1210
rect -5100 1190 -5090 1210
rect -5040 1190 -5030 1210
rect -5010 1190 -4940 1210
rect -4920 1190 -4910 1210
rect -4860 1190 -4850 1210
rect -4830 1190 -4760 1210
rect -4740 1190 -4730 1210
rect -4680 1190 -4670 1210
rect -4650 1190 -4580 1210
rect -4560 1190 -4550 1210
rect -4500 1190 -4490 1210
rect -4470 1190 -4400 1210
rect -4380 1190 -4370 1210
rect -4320 1190 -4310 1210
rect -4290 1190 -4220 1210
rect -4200 1190 -4190 1210
rect -4140 1190 -4130 1210
rect -4110 1190 -4040 1210
rect -4020 1190 -4010 1210
rect -3960 1190 -3950 1210
rect -3930 1190 -3860 1210
rect -3840 1190 -3830 1210
rect -3780 1190 -3770 1210
rect -3750 1190 -3680 1210
rect -3660 1190 -3650 1210
rect -3600 1190 -3590 1210
rect -3570 1190 -3500 1210
rect -3480 1190 -3470 1210
rect -3420 1190 -3410 1210
rect -3390 1190 -3320 1210
rect -3300 1190 -3290 1210
rect -3240 1190 -3230 1210
rect -3210 1190 -3140 1210
rect -3120 1190 -3110 1210
rect -3060 1190 -3050 1210
rect -3030 1190 -2960 1210
rect -2940 1190 -2930 1210
rect -2880 1190 -2870 1210
rect -2850 1190 -2780 1210
rect -2760 1190 -2750 1210
rect -2700 1190 -2690 1210
rect -2670 1190 -2600 1210
rect -2580 1190 -2570 1210
rect -2520 1190 -2510 1210
rect -2490 1190 -2420 1210
rect -2400 1190 -2390 1210
rect -2340 1190 -2330 1210
rect -2310 1190 -2240 1210
rect -2220 1190 -2210 1210
rect -2160 1190 -2150 1210
rect -2130 1190 -2060 1210
rect -2040 1190 -2030 1210
rect -1980 1190 -1970 1210
rect -1950 1190 -1880 1210
rect -1860 1190 -1850 1210
rect -1800 1190 -1790 1210
rect -1770 1190 -1700 1210
rect -1680 1190 -1670 1210
rect -1620 1190 -1610 1210
rect -1590 1190 -1520 1210
rect -1500 1190 -1490 1210
rect -1440 1190 -1430 1210
rect -1410 1190 -1340 1210
rect -1320 1190 -1310 1210
rect -1260 1190 -1250 1210
rect -1230 1190 -1160 1210
rect -1140 1190 -1130 1210
rect -1080 1190 -1070 1210
rect -1050 1190 -980 1210
rect -960 1190 -950 1210
rect -900 1190 -890 1210
rect -870 1190 -800 1210
rect -780 1190 -770 1210
rect -725 1190 -710 1210
rect -690 1190 -620 1210
rect -600 1190 -530 1210
rect -510 1190 -440 1210
rect -420 1190 -350 1210
rect -330 1190 -260 1210
rect -240 1190 -170 1210
rect -150 1190 -80 1210
rect -60 1190 -50 1210
rect -11555 1155 -11535 1165
rect -11555 1065 -11535 1075
rect -11465 1155 -11445 1165
rect -11465 1065 -11445 1075
rect -11375 1155 -11355 1165
rect -11375 1065 -11355 1075
rect -11285 1155 -11265 1190
rect -11285 1065 -11265 1075
rect -11195 1155 -11175 1165
rect -11195 1065 -11175 1075
rect -11105 1155 -11085 1190
rect -11105 1065 -11085 1075
rect -11015 1155 -10995 1165
rect -11015 1065 -10995 1075
rect -10925 1155 -10905 1165
rect -10925 1065 -10905 1075
rect -10835 1155 -10815 1165
rect -10835 1065 -10815 1075
rect -10745 1155 -10725 1165
rect -10745 1065 -10725 1075
rect -10655 1155 -10635 1165
rect -10655 1065 -10635 1075
rect -10565 1155 -10545 1165
rect -10565 1065 -10545 1075
rect -10475 1155 -10455 1165
rect -10475 1065 -10455 1075
rect -10385 1155 -10365 1165
rect -10385 1065 -10365 1075
rect -10295 1155 -10275 1165
rect -10295 1065 -10275 1075
rect -10205 1155 -10185 1165
rect -10205 1065 -10185 1075
rect -10115 1155 -10095 1165
rect -10115 1065 -10095 1075
rect -10025 1155 -10005 1165
rect -10025 1065 -10005 1075
rect -9935 1155 -9915 1165
rect -9935 1065 -9915 1075
rect -9845 1155 -9825 1165
rect -9845 1065 -9825 1075
rect -9755 1155 -9735 1165
rect -9755 1065 -9735 1075
rect -9665 1155 -9645 1165
rect -9665 1065 -9645 1075
rect -9575 1155 -9555 1165
rect -9575 1065 -9555 1075
rect -9485 1155 -9465 1165
rect -9485 1065 -9465 1075
rect -9395 1155 -9375 1165
rect -9395 1065 -9375 1075
rect -9305 1155 -9285 1165
rect -9305 1065 -9285 1075
rect -9215 1155 -9195 1165
rect -9215 1065 -9195 1075
rect -9125 1155 -9105 1165
rect -9125 1065 -9105 1075
rect -9035 1155 -9015 1165
rect -9035 1065 -9015 1075
rect -8945 1155 -8925 1165
rect -8945 1065 -8925 1075
rect -8855 1155 -8835 1165
rect -8855 1065 -8835 1075
rect -8765 1155 -8745 1165
rect -8765 1065 -8745 1075
rect -8675 1155 -8655 1165
rect -8675 1065 -8655 1075
rect -8585 1155 -8565 1165
rect -8585 1065 -8565 1075
rect -8495 1155 -8475 1165
rect -8495 1065 -8475 1075
rect -8405 1155 -8385 1165
rect -8405 1065 -8385 1075
rect -8315 1155 -8295 1165
rect -8315 1065 -8295 1075
rect -8225 1155 -8205 1165
rect -8225 1065 -8205 1075
rect -8135 1155 -8115 1165
rect -8135 1065 -8115 1075
rect -8045 1155 -8025 1165
rect -8045 1065 -8025 1075
rect -7955 1155 -7935 1165
rect -7955 1065 -7935 1075
rect -7865 1155 -7845 1165
rect -7865 1065 -7845 1075
rect -7775 1155 -7755 1165
rect -7775 1065 -7755 1075
rect -7685 1155 -7665 1165
rect -7685 1065 -7665 1075
rect -7595 1155 -7575 1165
rect -7595 1065 -7575 1075
rect -7505 1155 -7485 1165
rect -7505 1065 -7485 1075
rect -7415 1155 -7395 1165
rect -7415 1065 -7395 1075
rect -7325 1155 -7305 1165
rect -7325 1065 -7305 1075
rect -7235 1155 -7215 1165
rect -7235 1065 -7215 1075
rect -7145 1155 -7125 1165
rect -7145 1065 -7125 1075
rect -7055 1155 -7035 1165
rect -7055 1065 -7035 1075
rect -6965 1155 -6945 1165
rect -6965 1065 -6945 1075
rect -6875 1155 -6855 1165
rect -6875 1065 -6855 1075
rect -6785 1155 -6765 1165
rect -6785 1065 -6765 1075
rect -6695 1155 -6675 1165
rect -6695 1065 -6675 1075
rect -6605 1155 -6585 1165
rect -6605 1065 -6585 1075
rect -6515 1155 -6495 1165
rect -6515 1065 -6495 1075
rect -6425 1155 -6405 1165
rect -6425 1065 -6405 1075
rect -6335 1155 -6315 1165
rect -6335 1065 -6315 1075
rect -6245 1155 -6225 1165
rect -6245 1065 -6225 1075
rect -6155 1155 -6135 1165
rect -6155 1065 -6135 1075
rect -6065 1155 -6045 1165
rect -6065 1065 -6045 1075
rect -5975 1155 -5955 1165
rect -5975 1065 -5955 1075
rect -5885 1155 -5865 1165
rect -5885 1065 -5865 1075
rect -5795 1155 -5775 1165
rect -5795 1065 -5775 1075
rect -5705 1155 -5685 1165
rect -5705 1065 -5685 1075
rect -5615 1155 -5595 1165
rect -5615 1065 -5595 1075
rect -5525 1155 -5505 1165
rect -5525 1065 -5505 1075
rect -5435 1155 -5415 1165
rect -5435 1065 -5415 1075
rect -5345 1155 -5325 1165
rect -5345 1065 -5325 1075
rect -5255 1155 -5235 1165
rect -5255 1065 -5235 1075
rect -5165 1155 -5145 1165
rect -5165 1065 -5145 1075
rect -5075 1155 -5055 1165
rect -5075 1065 -5055 1075
rect -4985 1155 -4965 1165
rect -4985 1065 -4965 1075
rect -4895 1155 -4875 1165
rect -4895 1065 -4875 1075
rect -4805 1155 -4785 1165
rect -4805 1065 -4785 1075
rect -4715 1155 -4695 1165
rect -4715 1065 -4695 1075
rect -4625 1155 -4605 1165
rect -4625 1065 -4605 1075
rect -4535 1155 -4515 1165
rect -4535 1065 -4515 1075
rect -4445 1155 -4425 1165
rect -4445 1065 -4425 1075
rect -4355 1155 -4335 1165
rect -4355 1065 -4335 1075
rect -4265 1155 -4245 1165
rect -4265 1065 -4245 1075
rect -4175 1155 -4155 1165
rect -4175 1065 -4155 1075
rect -4085 1155 -4065 1165
rect -4085 1065 -4065 1075
rect -3995 1155 -3975 1165
rect -3995 1065 -3975 1075
rect -3905 1155 -3885 1165
rect -3905 1065 -3885 1075
rect -3815 1155 -3795 1165
rect -3815 1065 -3795 1075
rect -3725 1155 -3705 1165
rect -3725 1065 -3705 1075
rect -3635 1155 -3615 1165
rect -3635 1065 -3615 1075
rect -3545 1155 -3525 1165
rect -3545 1065 -3525 1075
rect -3455 1155 -3435 1165
rect -3455 1065 -3435 1075
rect -3365 1155 -3345 1165
rect -3365 1065 -3345 1075
rect -3275 1155 -3255 1165
rect -3275 1065 -3255 1075
rect -3185 1155 -3165 1165
rect -3185 1065 -3165 1075
rect -3095 1155 -3075 1165
rect -3095 1065 -3075 1075
rect -3005 1155 -2985 1165
rect -3005 1065 -2985 1075
rect -2915 1155 -2895 1165
rect -2915 1065 -2895 1075
rect -2825 1155 -2805 1165
rect -2825 1065 -2805 1075
rect -2735 1155 -2715 1165
rect -2735 1065 -2715 1075
rect -2645 1155 -2625 1165
rect -2645 1065 -2625 1075
rect -2555 1155 -2535 1165
rect -2555 1065 -2535 1075
rect -2465 1155 -2445 1165
rect -2465 1065 -2445 1075
rect -2375 1155 -2355 1165
rect -2375 1065 -2355 1075
rect -2285 1155 -2265 1165
rect -2285 1065 -2265 1075
rect -2195 1155 -2175 1165
rect -2195 1065 -2175 1075
rect -2105 1155 -2085 1165
rect -2105 1065 -2085 1075
rect -2015 1155 -1995 1165
rect -2015 1065 -1995 1075
rect -1925 1155 -1905 1165
rect -1925 1065 -1905 1075
rect -1835 1155 -1815 1165
rect -1835 1065 -1815 1075
rect -1745 1155 -1725 1165
rect -1745 1065 -1725 1075
rect -1655 1155 -1635 1165
rect -1655 1065 -1635 1075
rect -1565 1155 -1545 1165
rect -1565 1065 -1545 1075
rect -1475 1155 -1455 1165
rect -1475 1065 -1455 1075
rect -1385 1155 -1365 1165
rect -1385 1065 -1365 1075
rect -1295 1155 -1275 1165
rect -1295 1065 -1275 1075
rect -1205 1155 -1185 1165
rect -1205 1065 -1185 1075
rect -1115 1155 -1095 1165
rect -1115 1065 -1095 1075
rect -1025 1155 -1005 1165
rect -1025 1065 -1005 1075
rect -935 1155 -915 1165
rect -935 1065 -915 1075
rect -845 1155 -825 1165
rect -845 1065 -825 1075
rect -755 1155 -735 1165
rect -755 1065 -735 1075
rect -665 1155 -645 1165
rect -665 1065 -645 1075
rect -575 1155 -555 1165
rect -575 1065 -555 1075
rect -485 1155 -465 1190
rect -485 1065 -465 1075
rect -395 1155 -375 1165
rect -395 1065 -375 1075
rect -305 1155 -285 1190
rect -305 1065 -285 1075
rect -215 1155 -195 1165
rect -215 1065 -195 1075
rect -125 1155 -105 1165
rect -125 1065 -105 1075
rect -35 1155 -15 1165
rect -35 1065 -15 1075
rect 25 1035 45 1235
rect -11615 1015 -11555 1035
rect -11535 1015 -11510 1035
rect -11490 1015 -11420 1035
rect -11400 1015 -11330 1035
rect -11310 1015 -11240 1035
rect -11220 1015 -11150 1035
rect -11130 1015 -11060 1035
rect -11040 1015 -10970 1035
rect -10950 1015 -10880 1035
rect -10860 1015 -10835 1035
rect -10815 1015 -10790 1035
rect -10770 1015 -10700 1035
rect -10680 1015 -10655 1035
rect -10635 1015 -10610 1035
rect -10590 1015 -10520 1035
rect -10500 1015 -10475 1035
rect -10455 1015 -10430 1035
rect -10410 1015 -10340 1035
rect -10320 1015 -10295 1035
rect -10275 1015 -10250 1035
rect -10230 1015 -10160 1035
rect -10140 1015 -10115 1035
rect -10095 1015 -10070 1035
rect -10050 1015 -9980 1035
rect -9960 1015 -9935 1035
rect -9915 1015 -9890 1035
rect -9870 1015 -9800 1035
rect -9780 1015 -9755 1035
rect -9735 1015 -9710 1035
rect -9690 1015 -9620 1035
rect -9600 1015 -9575 1035
rect -9555 1015 -9530 1035
rect -9510 1015 -9440 1035
rect -9420 1015 -9395 1035
rect -9375 1015 -9350 1035
rect -9330 1015 -9260 1035
rect -9240 1015 -9215 1035
rect -9195 1015 -9170 1035
rect -9150 1015 -9080 1035
rect -9060 1015 -9035 1035
rect -9015 1015 -8990 1035
rect -8970 1015 -8900 1035
rect -8880 1015 -8855 1035
rect -8835 1015 -8810 1035
rect -8790 1015 -8720 1035
rect -8700 1015 -8675 1035
rect -8655 1015 -8630 1035
rect -8610 1015 -8540 1035
rect -8520 1015 -8495 1035
rect -8475 1015 -8450 1035
rect -8430 1015 -8360 1035
rect -8340 1015 -8315 1035
rect -8295 1015 -8270 1035
rect -8250 1015 -8180 1035
rect -8160 1015 -8135 1035
rect -8115 1015 -8090 1035
rect -8070 1015 -8000 1035
rect -7980 1015 -7955 1035
rect -7935 1015 -7910 1035
rect -7890 1015 -7820 1035
rect -7800 1015 -7775 1035
rect -7755 1015 -7730 1035
rect -7710 1015 -7640 1035
rect -7620 1015 -7595 1035
rect -7575 1015 -7550 1035
rect -7530 1015 -7460 1035
rect -7440 1015 -7415 1035
rect -7395 1015 -7370 1035
rect -7350 1015 -7280 1035
rect -7260 1015 -7235 1035
rect -7215 1015 -7190 1035
rect -7170 1015 -7100 1035
rect -7080 1015 -7055 1035
rect -7035 1015 -7010 1035
rect -6990 1015 -6920 1035
rect -6900 1015 -6875 1035
rect -6855 1015 -6830 1035
rect -6810 1015 -6740 1035
rect -6720 1015 -6695 1035
rect -6675 1015 -6650 1035
rect -6630 1015 -6560 1035
rect -6540 1015 -6515 1035
rect -6495 1015 -6470 1035
rect -6450 1015 -6380 1035
rect -6360 1015 -6335 1035
rect -6315 1015 -6290 1035
rect -6270 1015 -6200 1035
rect -6180 1015 -6155 1035
rect -6135 1015 -6110 1035
rect -6090 1015 -6020 1035
rect -6000 1015 -5975 1035
rect -5955 1015 -5930 1035
rect -5910 1015 -5840 1035
rect -5820 1015 -5795 1035
rect -5775 1015 -5750 1035
rect -5730 1015 -5660 1035
rect -5640 1015 -5615 1035
rect -5595 1015 -5570 1035
rect -5550 1015 -5480 1035
rect -5460 1015 -5435 1035
rect -5415 1015 -5390 1035
rect -5370 1015 -5300 1035
rect -5280 1015 -5255 1035
rect -5235 1015 -5210 1035
rect -5190 1015 -5120 1035
rect -5100 1015 -5075 1035
rect -5055 1015 -5030 1035
rect -5010 1015 -4940 1035
rect -4920 1015 -4895 1035
rect -4875 1015 -4850 1035
rect -4830 1015 -4760 1035
rect -4740 1015 -4715 1035
rect -4695 1015 -4670 1035
rect -4650 1015 -4580 1035
rect -4560 1015 -4535 1035
rect -4515 1015 -4490 1035
rect -4470 1015 -4400 1035
rect -4380 1015 -4355 1035
rect -4335 1015 -4310 1035
rect -4290 1015 -4220 1035
rect -4200 1015 -4175 1035
rect -4155 1015 -4130 1035
rect -4110 1015 -4040 1035
rect -4020 1015 -3995 1035
rect -3975 1015 -3950 1035
rect -3930 1015 -3860 1035
rect -3840 1015 -3815 1035
rect -3795 1015 -3770 1035
rect -3750 1015 -3680 1035
rect -3660 1015 -3635 1035
rect -3615 1015 -3590 1035
rect -3570 1015 -3500 1035
rect -3480 1015 -3455 1035
rect -3435 1015 -3410 1035
rect -3390 1015 -3320 1035
rect -3300 1015 -3275 1035
rect -3255 1015 -3230 1035
rect -3210 1015 -3140 1035
rect -3120 1015 -3095 1035
rect -3075 1015 -3050 1035
rect -3030 1015 -2960 1035
rect -2940 1015 -2915 1035
rect -2895 1015 -2870 1035
rect -2850 1015 -2780 1035
rect -2760 1015 -2735 1035
rect -2715 1015 -2690 1035
rect -2670 1015 -2600 1035
rect -2580 1015 -2555 1035
rect -2535 1015 -2510 1035
rect -2490 1015 -2420 1035
rect -2400 1015 -2375 1035
rect -2355 1015 -2330 1035
rect -2310 1015 -2240 1035
rect -2220 1015 -2195 1035
rect -2175 1015 -2150 1035
rect -2130 1015 -2060 1035
rect -2040 1015 -2015 1035
rect -1995 1015 -1970 1035
rect -1950 1015 -1880 1035
rect -1860 1015 -1835 1035
rect -1815 1015 -1790 1035
rect -1770 1015 -1700 1035
rect -1680 1015 -1655 1035
rect -1635 1015 -1610 1035
rect -1590 1015 -1520 1035
rect -1500 1015 -1475 1035
rect -1455 1015 -1430 1035
rect -1410 1015 -1340 1035
rect -1320 1015 -1295 1035
rect -1275 1015 -1250 1035
rect -1230 1015 -1160 1035
rect -1140 1015 -1115 1035
rect -1095 1015 -1070 1035
rect -1050 1015 -980 1035
rect -960 1015 -935 1035
rect -915 1015 -890 1035
rect -870 1015 -800 1035
rect -780 1015 -755 1035
rect -735 1015 -710 1035
rect -690 1015 -620 1035
rect -600 1015 -530 1035
rect -510 1015 -440 1035
rect -420 1015 -350 1035
rect -330 1015 -260 1035
rect -240 1015 -170 1035
rect -150 1015 -80 1035
rect -60 1015 -35 1035
rect -15 1015 45 1035
rect -11615 960 -11555 980
rect -11535 960 -11510 980
rect -11490 960 -11420 980
rect -11400 960 -11330 980
rect -11310 960 -11240 980
rect -11220 960 -11150 980
rect -11130 960 -11060 980
rect -11040 960 -10970 980
rect -10950 960 -10880 980
rect -10860 960 -10835 980
rect -10815 960 -10790 980
rect -10770 960 -10700 980
rect -10680 960 -10655 980
rect -10635 960 -10610 980
rect -10590 960 -10520 980
rect -10500 960 -10475 980
rect -10455 960 -10430 980
rect -10410 960 -10340 980
rect -10320 960 -10295 980
rect -10275 960 -10250 980
rect -10230 960 -10160 980
rect -10140 960 -10115 980
rect -10095 960 -10070 980
rect -10050 960 -9980 980
rect -9960 960 -9935 980
rect -9915 960 -9890 980
rect -9870 960 -9800 980
rect -9780 960 -9755 980
rect -9735 960 -9710 980
rect -9690 960 -9620 980
rect -9600 960 -9575 980
rect -9555 960 -9530 980
rect -9510 960 -9440 980
rect -9420 960 -9395 980
rect -9375 960 -9350 980
rect -9330 960 -9260 980
rect -9240 960 -9215 980
rect -9195 960 -9170 980
rect -9150 960 -9080 980
rect -9060 960 -9035 980
rect -9015 960 -8990 980
rect -8970 960 -8900 980
rect -8880 960 -8855 980
rect -8835 960 -8810 980
rect -8790 960 -8720 980
rect -8700 960 -8675 980
rect -8655 960 -8630 980
rect -8610 960 -8540 980
rect -8520 960 -8495 980
rect -8475 960 -8450 980
rect -8430 960 -8360 980
rect -8340 960 -8315 980
rect -8295 960 -8270 980
rect -8250 960 -8180 980
rect -8160 960 -8135 980
rect -8115 960 -8090 980
rect -8070 960 -8000 980
rect -7980 960 -7955 980
rect -7935 960 -7910 980
rect -7890 960 -7820 980
rect -7800 960 -7775 980
rect -7755 960 -7730 980
rect -7710 960 -7640 980
rect -7620 960 -7595 980
rect -7575 960 -7550 980
rect -7530 960 -7460 980
rect -7440 960 -7415 980
rect -7395 960 -7370 980
rect -7350 960 -7280 980
rect -7260 960 -7235 980
rect -7215 960 -7190 980
rect -7170 960 -7100 980
rect -7080 960 -7055 980
rect -7035 960 -7010 980
rect -6990 960 -6920 980
rect -6900 960 -6875 980
rect -6855 960 -6830 980
rect -6810 960 -6740 980
rect -6720 960 -6695 980
rect -6675 960 -6650 980
rect -6630 960 -6560 980
rect -6540 960 -6515 980
rect -6495 960 -6470 980
rect -6450 960 -6380 980
rect -6360 960 -6335 980
rect -6315 960 -6290 980
rect -6270 960 -6200 980
rect -6180 960 -6155 980
rect -6135 960 -6110 980
rect -6090 960 -6020 980
rect -6000 960 -5975 980
rect -5955 960 -5930 980
rect -5910 960 -5840 980
rect -5820 960 -5795 980
rect -5775 960 -5750 980
rect -5730 960 -5660 980
rect -5640 960 -5615 980
rect -5595 960 -5570 980
rect -5550 960 -5480 980
rect -5460 960 -5435 980
rect -5415 960 -5390 980
rect -5370 960 -5300 980
rect -5280 960 -5255 980
rect -5235 960 -5210 980
rect -5190 960 -5120 980
rect -5100 960 -5075 980
rect -5055 960 -5030 980
rect -5010 960 -4940 980
rect -4920 960 -4895 980
rect -4875 960 -4850 980
rect -4830 960 -4760 980
rect -4740 960 -4715 980
rect -4695 960 -4670 980
rect -4650 960 -4580 980
rect -4560 960 -4535 980
rect -4515 960 -4490 980
rect -4470 960 -4400 980
rect -4380 960 -4355 980
rect -4335 960 -4310 980
rect -4290 960 -4220 980
rect -4200 960 -4175 980
rect -4155 960 -4130 980
rect -4110 960 -4040 980
rect -4020 960 -3995 980
rect -3975 960 -3950 980
rect -3930 960 -3860 980
rect -3840 960 -3815 980
rect -3795 960 -3770 980
rect -3750 960 -3680 980
rect -3660 960 -3635 980
rect -3615 960 -3590 980
rect -3570 960 -3500 980
rect -3480 960 -3455 980
rect -3435 960 -3410 980
rect -3390 960 -3320 980
rect -3300 960 -3275 980
rect -3255 960 -3230 980
rect -3210 960 -3140 980
rect -3120 960 -3095 980
rect -3075 960 -3050 980
rect -3030 960 -2960 980
rect -2940 960 -2915 980
rect -2895 960 -2870 980
rect -2850 960 -2780 980
rect -2760 960 -2735 980
rect -2715 960 -2690 980
rect -2670 960 -2600 980
rect -2580 960 -2555 980
rect -2535 960 -2510 980
rect -2490 960 -2420 980
rect -2400 960 -2375 980
rect -2355 960 -2330 980
rect -2310 960 -2240 980
rect -2220 960 -2195 980
rect -2175 960 -2150 980
rect -2130 960 -2060 980
rect -2040 960 -2015 980
rect -1995 960 -1970 980
rect -1950 960 -1880 980
rect -1860 960 -1835 980
rect -1815 960 -1790 980
rect -1770 960 -1700 980
rect -1680 960 -1655 980
rect -1635 960 -1610 980
rect -1590 960 -1520 980
rect -1500 960 -1475 980
rect -1455 960 -1430 980
rect -1410 960 -1340 980
rect -1320 960 -1295 980
rect -1275 960 -1250 980
rect -1230 960 -1160 980
rect -1140 960 -1115 980
rect -1095 960 -1070 980
rect -1050 960 -980 980
rect -960 960 -935 980
rect -915 960 -890 980
rect -870 960 -800 980
rect -780 960 -755 980
rect -735 960 -710 980
rect -690 960 -620 980
rect -600 960 -530 980
rect -510 960 -440 980
rect -420 960 -350 980
rect -330 960 -260 980
rect -240 960 -170 980
rect -150 960 -80 980
rect -60 960 -35 980
rect -15 960 45 980
rect -11615 760 -11595 960
rect -11555 920 -11535 930
rect -11555 830 -11535 840
rect -11465 920 -11445 930
rect -11465 830 -11445 840
rect -11375 920 -11355 930
rect -11375 830 -11355 840
rect -11285 920 -11265 930
rect -11285 805 -11265 840
rect -11195 920 -11175 930
rect -11195 830 -11175 840
rect -11105 920 -11085 930
rect -11105 805 -11085 840
rect -11015 920 -10995 930
rect -11015 830 -10995 840
rect -10925 920 -10905 930
rect -10925 830 -10905 840
rect -10835 920 -10815 930
rect -10835 830 -10815 840
rect -10745 920 -10725 930
rect -10745 830 -10725 840
rect -10655 920 -10635 930
rect -10655 830 -10635 840
rect -10565 920 -10545 930
rect -10565 830 -10545 840
rect -10475 920 -10455 930
rect -10475 830 -10455 840
rect -10385 920 -10365 930
rect -10385 830 -10365 840
rect -10295 920 -10275 930
rect -10295 830 -10275 840
rect -10205 920 -10185 930
rect -10205 830 -10185 840
rect -10115 920 -10095 930
rect -10115 830 -10095 840
rect -10025 920 -10005 930
rect -10025 830 -10005 840
rect -9935 920 -9915 930
rect -9935 830 -9915 840
rect -9845 920 -9825 930
rect -9845 830 -9825 840
rect -9755 920 -9735 930
rect -9755 830 -9735 840
rect -9665 920 -9645 930
rect -9665 830 -9645 840
rect -9575 920 -9555 930
rect -9575 830 -9555 840
rect -9485 920 -9465 930
rect -9485 830 -9465 840
rect -9395 920 -9375 930
rect -9395 830 -9375 840
rect -9305 920 -9285 930
rect -9305 830 -9285 840
rect -9215 920 -9195 930
rect -9215 830 -9195 840
rect -9125 920 -9105 930
rect -9125 830 -9105 840
rect -9035 920 -9015 930
rect -9035 830 -9015 840
rect -8945 920 -8925 930
rect -8945 830 -8925 840
rect -8855 920 -8835 930
rect -8855 830 -8835 840
rect -8765 920 -8745 930
rect -8765 830 -8745 840
rect -8675 920 -8655 930
rect -8675 830 -8655 840
rect -8585 920 -8565 930
rect -8585 830 -8565 840
rect -8495 920 -8475 930
rect -8495 830 -8475 840
rect -8405 920 -8385 930
rect -8405 830 -8385 840
rect -8315 920 -8295 930
rect -8315 830 -8295 840
rect -8225 920 -8205 930
rect -8225 830 -8205 840
rect -8135 920 -8115 930
rect -8135 830 -8115 840
rect -8045 920 -8025 930
rect -8045 830 -8025 840
rect -7955 920 -7935 930
rect -7955 830 -7935 840
rect -7865 920 -7845 930
rect -7865 830 -7845 840
rect -7775 920 -7755 930
rect -7775 830 -7755 840
rect -7685 920 -7665 930
rect -7685 830 -7665 840
rect -7595 920 -7575 930
rect -7595 830 -7575 840
rect -7505 920 -7485 930
rect -7505 830 -7485 840
rect -7415 920 -7395 930
rect -7415 830 -7395 840
rect -7325 920 -7305 930
rect -7325 830 -7305 840
rect -7235 920 -7215 930
rect -7235 830 -7215 840
rect -7145 920 -7125 930
rect -7145 830 -7125 840
rect -7055 920 -7035 930
rect -7055 830 -7035 840
rect -6965 920 -6945 930
rect -6965 830 -6945 840
rect -6875 920 -6855 930
rect -6875 830 -6855 840
rect -6785 920 -6765 930
rect -6785 830 -6765 840
rect -6695 920 -6675 930
rect -6695 830 -6675 840
rect -6605 920 -6585 930
rect -6605 830 -6585 840
rect -6515 920 -6495 930
rect -6515 830 -6495 840
rect -6425 920 -6405 930
rect -6425 830 -6405 840
rect -6335 920 -6315 930
rect -6335 830 -6315 840
rect -6245 920 -6225 930
rect -6245 830 -6225 840
rect -6155 920 -6135 930
rect -6155 830 -6135 840
rect -6065 920 -6045 930
rect -6065 830 -6045 840
rect -5975 920 -5955 930
rect -5975 830 -5955 840
rect -5885 920 -5865 930
rect -5885 830 -5865 840
rect -5795 920 -5775 930
rect -5795 830 -5775 840
rect -5705 920 -5685 930
rect -5705 830 -5685 840
rect -5615 920 -5595 930
rect -5615 830 -5595 840
rect -5525 920 -5505 930
rect -5525 830 -5505 840
rect -5435 920 -5415 930
rect -5435 830 -5415 840
rect -5345 920 -5325 930
rect -5345 830 -5325 840
rect -5255 920 -5235 930
rect -5255 830 -5235 840
rect -5165 920 -5145 930
rect -5165 830 -5145 840
rect -5075 920 -5055 930
rect -5075 830 -5055 840
rect -4985 920 -4965 930
rect -4985 830 -4965 840
rect -4895 920 -4875 930
rect -4895 830 -4875 840
rect -4805 920 -4785 930
rect -4805 830 -4785 840
rect -4715 920 -4695 930
rect -4715 830 -4695 840
rect -4625 920 -4605 930
rect -4625 830 -4605 840
rect -4535 920 -4515 930
rect -4535 830 -4515 840
rect -4445 920 -4425 930
rect -4445 830 -4425 840
rect -4355 920 -4335 930
rect -4355 830 -4335 840
rect -4265 920 -4245 930
rect -4265 830 -4245 840
rect -4175 920 -4155 930
rect -4175 830 -4155 840
rect -4085 920 -4065 930
rect -4085 830 -4065 840
rect -3995 920 -3975 930
rect -3995 830 -3975 840
rect -3905 920 -3885 930
rect -3905 830 -3885 840
rect -3815 920 -3795 930
rect -3815 830 -3795 840
rect -3725 920 -3705 930
rect -3725 830 -3705 840
rect -3635 920 -3615 930
rect -3635 830 -3615 840
rect -3545 920 -3525 930
rect -3545 830 -3525 840
rect -3455 920 -3435 930
rect -3455 830 -3435 840
rect -3365 920 -3345 930
rect -3365 830 -3345 840
rect -3275 920 -3255 930
rect -3275 830 -3255 840
rect -3185 920 -3165 930
rect -3185 830 -3165 840
rect -3095 920 -3075 930
rect -3095 830 -3075 840
rect -3005 920 -2985 930
rect -3005 830 -2985 840
rect -2915 920 -2895 930
rect -2915 830 -2895 840
rect -2825 920 -2805 930
rect -2825 830 -2805 840
rect -2735 920 -2715 930
rect -2735 830 -2715 840
rect -2645 920 -2625 930
rect -2645 830 -2625 840
rect -2555 920 -2535 930
rect -2555 830 -2535 840
rect -2465 920 -2445 930
rect -2465 830 -2445 840
rect -2375 920 -2355 930
rect -2375 830 -2355 840
rect -2285 920 -2265 930
rect -2285 830 -2265 840
rect -2195 920 -2175 930
rect -2195 830 -2175 840
rect -2105 920 -2085 930
rect -2105 830 -2085 840
rect -2015 920 -1995 930
rect -2015 830 -1995 840
rect -1925 920 -1905 930
rect -1925 830 -1905 840
rect -1835 920 -1815 930
rect -1835 830 -1815 840
rect -1745 920 -1725 930
rect -1745 830 -1725 840
rect -1655 920 -1635 930
rect -1655 830 -1635 840
rect -1565 920 -1545 930
rect -1565 830 -1545 840
rect -1475 920 -1455 930
rect -1475 830 -1455 840
rect -1385 920 -1365 930
rect -1385 830 -1365 840
rect -1295 920 -1275 930
rect -1295 830 -1275 840
rect -1205 920 -1185 930
rect -1205 830 -1185 840
rect -1115 920 -1095 930
rect -1115 830 -1095 840
rect -1025 920 -1005 930
rect -1025 830 -1005 840
rect -935 920 -915 930
rect -935 830 -915 840
rect -845 920 -825 930
rect -845 830 -825 840
rect -755 920 -735 930
rect -755 830 -735 840
rect -665 920 -645 930
rect -665 830 -645 840
rect -575 920 -555 930
rect -575 830 -555 840
rect -485 920 -465 930
rect -485 805 -465 840
rect -395 920 -375 930
rect -395 830 -375 840
rect -305 920 -285 930
rect -305 805 -285 840
rect -215 920 -195 930
rect -215 830 -195 840
rect -125 920 -105 930
rect -125 830 -105 840
rect -35 920 -15 930
rect -35 830 -15 840
rect -11520 785 -11510 805
rect -11490 785 -11420 805
rect -11400 785 -11330 805
rect -11310 785 -11240 805
rect -11220 785 -11150 805
rect -11130 785 -11060 805
rect -11040 785 -10970 805
rect -10950 785 -10880 805
rect -10860 785 -10845 805
rect -10800 785 -10790 805
rect -10770 785 -10700 805
rect -10680 785 -10670 805
rect -10620 785 -10610 805
rect -10590 785 -10520 805
rect -10500 785 -10490 805
rect -10440 785 -10430 805
rect -10410 785 -10340 805
rect -10320 785 -10310 805
rect -10260 785 -10250 805
rect -10230 785 -10160 805
rect -10140 785 -10130 805
rect -10080 785 -10070 805
rect -10050 785 -9980 805
rect -9960 785 -9950 805
rect -9900 785 -9890 805
rect -9870 785 -9800 805
rect -9780 785 -9770 805
rect -9720 785 -9710 805
rect -9690 785 -9620 805
rect -9600 785 -9590 805
rect -9540 785 -9530 805
rect -9510 785 -9440 805
rect -9420 785 -9410 805
rect -9360 785 -9350 805
rect -9330 785 -9260 805
rect -9240 785 -9230 805
rect -9180 785 -9170 805
rect -9150 785 -9080 805
rect -9060 785 -9050 805
rect -9000 785 -8990 805
rect -8970 785 -8900 805
rect -8880 785 -8870 805
rect -8820 785 -8810 805
rect -8790 785 -8720 805
rect -8700 785 -8690 805
rect -8640 785 -8630 805
rect -8610 785 -8540 805
rect -8520 785 -8510 805
rect -8460 785 -8450 805
rect -8430 785 -8360 805
rect -8340 785 -8330 805
rect -8280 785 -8270 805
rect -8250 785 -8180 805
rect -8160 785 -8150 805
rect -8100 785 -8090 805
rect -8070 785 -8000 805
rect -7980 785 -7970 805
rect -7920 785 -7910 805
rect -7890 785 -7820 805
rect -7800 785 -7790 805
rect -7740 785 -7730 805
rect -7710 785 -7640 805
rect -7620 785 -7610 805
rect -7560 785 -7550 805
rect -7530 785 -7460 805
rect -7440 785 -7430 805
rect -7380 785 -7370 805
rect -7350 785 -7280 805
rect -7260 785 -7250 805
rect -7200 785 -7190 805
rect -7170 785 -7100 805
rect -7080 785 -7070 805
rect -7020 785 -7010 805
rect -6990 785 -6920 805
rect -6900 785 -6890 805
rect -6840 785 -6830 805
rect -6810 785 -6740 805
rect -6720 785 -6710 805
rect -6660 785 -6650 805
rect -6630 785 -6560 805
rect -6540 785 -6530 805
rect -6480 785 -6470 805
rect -6450 785 -6380 805
rect -6360 785 -6350 805
rect -6300 785 -6290 805
rect -6270 785 -6200 805
rect -6180 785 -6170 805
rect -6120 785 -6110 805
rect -6090 785 -6020 805
rect -6000 785 -5990 805
rect -5940 785 -5930 805
rect -5910 785 -5840 805
rect -5820 785 -5810 805
rect -5760 785 -5750 805
rect -5730 785 -5660 805
rect -5640 785 -5630 805
rect -5580 785 -5570 805
rect -5550 785 -5480 805
rect -5460 785 -5450 805
rect -5400 785 -5390 805
rect -5370 785 -5300 805
rect -5280 785 -5270 805
rect -5220 785 -5210 805
rect -5190 785 -5120 805
rect -5100 785 -5090 805
rect -5040 785 -5030 805
rect -5010 785 -4940 805
rect -4920 785 -4910 805
rect -4860 785 -4850 805
rect -4830 785 -4760 805
rect -4740 785 -4730 805
rect -4680 785 -4670 805
rect -4650 785 -4580 805
rect -4560 785 -4550 805
rect -4500 785 -4490 805
rect -4470 785 -4400 805
rect -4380 785 -4370 805
rect -4320 785 -4310 805
rect -4290 785 -4220 805
rect -4200 785 -4190 805
rect -4140 785 -4130 805
rect -4110 785 -4040 805
rect -4020 785 -4010 805
rect -3960 785 -3950 805
rect -3930 785 -3860 805
rect -3840 785 -3830 805
rect -3780 785 -3770 805
rect -3750 785 -3680 805
rect -3660 785 -3650 805
rect -3600 785 -3590 805
rect -3570 785 -3500 805
rect -3480 785 -3470 805
rect -3420 785 -3410 805
rect -3390 785 -3320 805
rect -3300 785 -3290 805
rect -3240 785 -3230 805
rect -3210 785 -3140 805
rect -3120 785 -3110 805
rect -3060 785 -3050 805
rect -3030 785 -2960 805
rect -2940 785 -2930 805
rect -2880 785 -2870 805
rect -2850 785 -2780 805
rect -2760 785 -2750 805
rect -2700 785 -2690 805
rect -2670 785 -2600 805
rect -2580 785 -2570 805
rect -2520 785 -2510 805
rect -2490 785 -2420 805
rect -2400 785 -2390 805
rect -2340 785 -2330 805
rect -2310 785 -2240 805
rect -2220 785 -2210 805
rect -2160 785 -2150 805
rect -2130 785 -2060 805
rect -2040 785 -2030 805
rect -1980 785 -1970 805
rect -1950 785 -1880 805
rect -1860 785 -1850 805
rect -1800 785 -1790 805
rect -1770 785 -1700 805
rect -1680 785 -1670 805
rect -1620 785 -1610 805
rect -1590 785 -1520 805
rect -1500 785 -1490 805
rect -1440 785 -1430 805
rect -1410 785 -1340 805
rect -1320 785 -1310 805
rect -1260 785 -1250 805
rect -1230 785 -1160 805
rect -1140 785 -1130 805
rect -1080 785 -1070 805
rect -1050 785 -980 805
rect -960 785 -950 805
rect -900 785 -890 805
rect -870 785 -800 805
rect -780 785 -770 805
rect -725 785 -710 805
rect -690 785 -620 805
rect -600 785 -530 805
rect -510 785 -440 805
rect -420 785 -350 805
rect -330 785 -260 805
rect -240 785 -170 805
rect -150 785 -80 805
rect -60 785 -50 805
rect 25 760 45 960
rect -11615 740 -11510 760
rect -11490 740 -11420 760
rect -11400 740 -11330 760
rect -11310 740 -11240 760
rect -11220 740 -11150 760
rect -11130 740 -11060 760
rect -11040 740 -10970 760
rect -10950 740 -10880 760
rect -10860 740 -10790 760
rect -10770 740 -10700 760
rect -10680 740 -10610 760
rect -10590 740 -10520 760
rect -10500 740 -10430 760
rect -10410 740 -10340 760
rect -10320 740 -10250 760
rect -10230 740 -10160 760
rect -10140 740 -10070 760
rect -10050 740 -9980 760
rect -9960 740 -9890 760
rect -9870 740 -9800 760
rect -9780 740 -9710 760
rect -9690 740 -9620 760
rect -9600 740 -9530 760
rect -9510 740 -9440 760
rect -9420 740 -9350 760
rect -9330 740 -9260 760
rect -9240 740 -9170 760
rect -9150 740 -9080 760
rect -9060 740 -8990 760
rect -8970 740 -8900 760
rect -8880 740 -8810 760
rect -8790 740 -8720 760
rect -8700 740 -8630 760
rect -8610 740 -8540 760
rect -8520 740 -8450 760
rect -8430 740 -8360 760
rect -8340 740 -8270 760
rect -8250 740 -8180 760
rect -8160 740 -8090 760
rect -8070 740 -8000 760
rect -7980 740 -7910 760
rect -7890 740 -7820 760
rect -7800 740 -7730 760
rect -7710 740 -7640 760
rect -7620 740 -7550 760
rect -7530 740 -7460 760
rect -7440 740 -7370 760
rect -7350 740 -7280 760
rect -7260 740 -7190 760
rect -7170 740 -7100 760
rect -7080 740 -7010 760
rect -6990 740 -6920 760
rect -6900 740 -6830 760
rect -6810 740 -6740 760
rect -6720 740 -6650 760
rect -6630 740 -6560 760
rect -6540 740 -6470 760
rect -6450 740 -6380 760
rect -6360 740 -6290 760
rect -6270 740 -6200 760
rect -6180 740 -6110 760
rect -6090 740 -6020 760
rect -6000 740 -5930 760
rect -5910 740 -5840 760
rect -5820 740 -5750 760
rect -5730 740 -5660 760
rect -5640 740 -5570 760
rect -5550 740 -5480 760
rect -5460 740 -5390 760
rect -5370 740 -5300 760
rect -5280 740 -5210 760
rect -5190 740 -5120 760
rect -5100 740 -5030 760
rect -5010 740 -4940 760
rect -4920 740 -4850 760
rect -4830 740 -4760 760
rect -4740 740 -4670 760
rect -4650 740 -4580 760
rect -4560 740 -4490 760
rect -4470 740 -4400 760
rect -4380 740 -4310 760
rect -4290 740 -4220 760
rect -4200 740 -4130 760
rect -4110 740 -4040 760
rect -4020 740 -3950 760
rect -3930 740 -3860 760
rect -3840 740 -3770 760
rect -3750 740 -3680 760
rect -3660 740 -3590 760
rect -3570 740 -3500 760
rect -3480 740 -3410 760
rect -3390 740 -3320 760
rect -3300 740 -3230 760
rect -3210 740 -3140 760
rect -3120 740 -3050 760
rect -3030 740 -2960 760
rect -2940 740 -2870 760
rect -2850 740 -2780 760
rect -2760 740 -2690 760
rect -2670 740 -2600 760
rect -2580 740 -2510 760
rect -2490 740 -2420 760
rect -2400 740 -2330 760
rect -2310 740 -2240 760
rect -2220 740 -2150 760
rect -2130 740 -2060 760
rect -2040 740 -1970 760
rect -1950 740 -1880 760
rect -1860 740 -1790 760
rect -1770 740 -1700 760
rect -1680 740 -1610 760
rect -1590 740 -1520 760
rect -1500 740 -1430 760
rect -1410 740 -1340 760
rect -1320 740 -1250 760
rect -1230 740 -1160 760
rect -1140 740 -1070 760
rect -1050 740 -980 760
rect -960 740 -890 760
rect -870 740 -800 760
rect -780 740 -710 760
rect -690 740 -620 760
rect -600 740 -530 760
rect -510 740 -440 760
rect -420 740 -350 760
rect -330 740 -260 760
rect -240 740 -170 760
rect -150 740 -80 760
rect -60 740 45 760
rect -11565 700 -10115 720
rect -10095 700 -9935 720
rect -9915 700 -9755 720
rect -9735 700 -9575 720
rect -9555 700 -9395 720
rect -9375 700 -9215 720
rect -9195 700 -9035 720
rect -9015 700 -8855 720
rect -8835 700 -8675 720
rect -8655 700 -8495 720
rect -8475 700 -8315 720
rect -8295 700 -8135 720
rect -8115 700 -7955 720
rect -7935 700 -6515 720
rect -6495 700 -6335 720
rect -6315 700 -6155 720
rect -6135 700 -5975 720
rect -5955 700 -5795 720
rect -5775 700 -5615 720
rect -5595 700 -5435 720
rect -5415 700 -5255 720
rect -5235 700 -5075 720
rect -5055 700 -4895 720
rect -4875 700 -4715 720
rect -4695 700 -4535 720
rect -4515 700 -4355 720
rect -4335 700 -575 720
rect -555 700 -5 720
rect 100 680 120 1315
rect -11690 660 -11510 680
rect -11490 660 -11420 680
rect -11400 660 -11330 680
rect -11310 660 -11240 680
rect -11220 660 -11150 680
rect -11130 660 -11060 680
rect -11040 660 -10970 680
rect -10950 660 -10880 680
rect -10860 660 -10790 680
rect -10770 660 -10700 680
rect -10680 660 -10610 680
rect -10590 660 -10520 680
rect -10500 660 -10430 680
rect -10410 660 -10340 680
rect -10320 660 -10250 680
rect -10230 660 -10160 680
rect -10140 660 -10070 680
rect -10050 660 -9980 680
rect -9960 660 -9890 680
rect -9870 660 -9800 680
rect -9780 660 -9710 680
rect -9690 660 -9620 680
rect -9600 660 -9530 680
rect -9510 660 -9440 680
rect -9420 660 -9350 680
rect -9330 660 -9260 680
rect -9240 660 -9170 680
rect -9150 660 -9080 680
rect -9060 660 -8990 680
rect -8970 660 -8900 680
rect -8880 660 -8810 680
rect -8790 660 -8720 680
rect -8700 660 -8630 680
rect -8610 660 -8540 680
rect -8520 660 -8450 680
rect -8430 660 -8360 680
rect -8340 660 -8270 680
rect -8250 660 -8180 680
rect -8160 660 -8090 680
rect -8070 660 -8000 680
rect -7980 660 -7910 680
rect -7890 660 -7820 680
rect -7800 660 -7730 680
rect -7710 660 -7640 680
rect -7620 660 -7550 680
rect -7530 660 -7460 680
rect -7440 660 -7370 680
rect -7350 660 -7280 680
rect -7260 660 -7190 680
rect -7170 660 -7100 680
rect -7080 660 -7010 680
rect -6990 660 -6920 680
rect -6900 660 -6830 680
rect -6810 660 -6740 680
rect -6720 660 -6650 680
rect -6630 660 -6560 680
rect -6540 660 -6470 680
rect -6450 660 -6380 680
rect -6360 660 -6290 680
rect -6270 660 -6200 680
rect -6180 660 -6110 680
rect -6090 660 -6020 680
rect -6000 660 -5930 680
rect -5910 660 -5840 680
rect -5820 660 -5750 680
rect -5730 660 -5660 680
rect -5640 660 -5570 680
rect -5550 660 -5480 680
rect -5460 660 -5390 680
rect -5370 660 -5300 680
rect -5280 660 -5210 680
rect -5190 660 -5120 680
rect -5100 660 -5030 680
rect -5010 660 -4940 680
rect -4920 660 -4850 680
rect -4830 660 -4760 680
rect -4740 660 -4670 680
rect -4650 660 -4580 680
rect -4560 660 -4490 680
rect -4470 660 -4400 680
rect -4380 660 -4310 680
rect -4290 660 -4220 680
rect -4200 660 -4130 680
rect -4110 660 -4040 680
rect -4020 660 -3950 680
rect -3930 660 -3860 680
rect -3840 660 -3770 680
rect -3750 660 -3680 680
rect -3660 660 -3590 680
rect -3570 660 -3500 680
rect -3480 660 -3410 680
rect -3390 660 -3320 680
rect -3300 660 -3230 680
rect -3210 660 -3140 680
rect -3120 660 -3050 680
rect -3030 660 -2960 680
rect -2940 660 -2870 680
rect -2850 660 -2780 680
rect -2760 660 -2690 680
rect -2670 660 -2600 680
rect -2580 660 -2510 680
rect -2490 660 -2420 680
rect -2400 660 -2330 680
rect -2310 660 -2240 680
rect -2220 660 -2150 680
rect -2130 660 -2060 680
rect -2040 660 -1970 680
rect -1950 660 -1880 680
rect -1860 660 -1790 680
rect -1770 660 -1700 680
rect -1680 660 -1610 680
rect -1590 660 -1520 680
rect -1500 660 -1430 680
rect -1410 660 -1340 680
rect -1320 660 -1250 680
rect -1230 660 -1160 680
rect -1140 660 -1070 680
rect -1050 660 -980 680
rect -960 660 -890 680
rect -870 660 -800 680
rect -780 660 -710 680
rect -690 660 -620 680
rect -600 660 -530 680
rect -510 660 -440 680
rect -420 660 -350 680
rect -330 660 -260 680
rect -240 660 -170 680
rect -150 660 -80 680
rect -60 660 120 680
rect -11565 620 -10700 640
rect -10680 620 -10520 640
rect -10500 620 -7460 640
rect -7440 620 -7280 640
rect -7260 620 -7100 640
rect -7080 620 -6920 640
rect -6900 620 -3860 640
rect -3840 620 -3680 640
rect -3660 620 -395 640
rect -375 620 -5 640
rect -11565 580 -10340 600
rect -10320 580 -10160 600
rect -10140 580 -7820 600
rect -7800 580 -7640 600
rect -7620 580 -6740 600
rect -6720 580 -6560 600
rect -6540 580 -4220 600
rect -4200 580 -4040 600
rect -4020 580 -3140 600
rect -3120 580 -2960 600
rect -2940 580 -2780 600
rect -2760 580 -2600 600
rect -2580 580 -1700 600
rect -1680 580 -1520 600
rect -1500 580 -1340 600
rect -1320 580 -1160 600
rect -1140 580 -305 600
rect -285 580 -5 600
rect -11565 540 -10115 560
rect -10095 540 -7955 560
rect -7935 540 -3500 560
rect -3480 540 -3320 560
rect -3300 540 -2915 560
rect -2895 540 -2420 560
rect -2400 540 -2240 560
rect -2220 540 -2060 560
rect -2040 540 -1880 560
rect -1860 540 -980 560
rect -960 540 -800 560
rect -780 540 -485 560
rect -465 540 -5 560
rect -11565 500 -11465 520
rect -11445 500 -6515 520
rect -6495 500 -4355 520
rect -4335 500 -1475 520
rect -1455 500 -5 520
rect -11565 460 -11375 480
rect -11355 460 -6380 480
rect -6360 460 -6200 480
rect -6180 460 -6020 480
rect -6000 460 -5840 480
rect -5820 460 -5660 480
rect -5640 460 -5480 480
rect -5460 460 -5300 480
rect -5280 460 -5120 480
rect -5100 460 -4940 480
rect -4920 460 -4760 480
rect -4740 460 -4580 480
rect -4560 460 -4400 480
rect -4380 460 -5 480
rect -11565 420 -11285 440
rect -11265 420 -9980 440
rect -9960 420 -9800 440
rect -9780 420 -9620 440
rect -9600 420 -9440 440
rect -9420 420 -9260 440
rect -9240 420 -9080 440
rect -9060 420 -8900 440
rect -8880 420 -8720 440
rect -8700 420 -8540 440
rect -8520 420 -8360 440
rect -8340 420 -8180 440
rect -8160 420 -8000 440
rect -7980 420 -5 440
rect -11565 380 -11195 400
rect -11175 380 -6875 400
rect -6855 380 -6425 400
rect -6405 380 -6245 400
rect -6225 380 -6065 400
rect -6045 380 -5885 400
rect -5865 380 -5705 400
rect -5685 380 -5525 400
rect -5505 380 -5345 400
rect -5325 380 -5165 400
rect -5145 380 -4985 400
rect -4965 380 -4805 400
rect -4785 380 -4625 400
rect -4605 380 -4445 400
rect -4425 380 -3995 400
rect -3975 380 -1835 400
rect -1815 380 -1115 400
rect -1095 380 -5 400
rect -11565 340 -11105 360
rect -11085 340 -10475 360
rect -10455 340 -10025 360
rect -10005 340 -9845 360
rect -9825 340 -9665 360
rect -9645 340 -9485 360
rect -9465 340 -9305 360
rect -9285 340 -9125 360
rect -9105 340 -8945 360
rect -8925 340 -8765 360
rect -8745 340 -8585 360
rect -8565 340 -8405 360
rect -8385 340 -8225 360
rect -8205 340 -8045 360
rect -8025 340 -7595 360
rect -7575 340 -3275 360
rect -3255 340 -2555 360
rect -2535 340 -5 360
rect -11565 300 -10430 320
rect -10410 300 -10250 320
rect -10230 300 -7910 320
rect -7890 300 -7730 320
rect -7710 300 -6830 320
rect -6810 300 -6650 320
rect -6630 300 -4310 320
rect -4290 300 -4130 320
rect -4110 300 -3230 320
rect -3210 300 -3050 320
rect -3030 300 -2870 320
rect -2850 300 -2690 320
rect -2670 300 -1790 320
rect -1770 300 -1610 320
rect -1590 300 -1430 320
rect -1410 300 -1250 320
rect -1230 300 -215 320
rect -195 300 -5 320
rect -11565 260 -10790 280
rect -10770 260 -10610 280
rect -10590 260 -7550 280
rect -7530 260 -7370 280
rect -7350 260 -7190 280
rect -7170 260 -7010 280
rect -6990 260 -3950 280
rect -3930 260 -3770 280
rect -3750 260 -3590 280
rect -3570 260 -3410 280
rect -3390 260 -2510 280
rect -2490 260 -2330 280
rect -2310 260 -2150 280
rect -2130 260 -1970 280
rect -1950 260 -1070 280
rect -1050 260 -890 280
rect -870 260 -125 280
rect -105 260 -5 280
rect -11690 220 -11510 240
rect -11490 220 -11420 240
rect -11400 220 -11330 240
rect -11310 220 -11240 240
rect -11220 220 -11150 240
rect -11130 220 -11060 240
rect -11040 220 -10970 240
rect -10950 220 -10880 240
rect -10860 220 -10790 240
rect -10770 220 -10700 240
rect -10680 220 -10610 240
rect -10590 220 -10520 240
rect -10500 220 -10430 240
rect -10410 220 -10340 240
rect -10320 220 -10250 240
rect -10230 220 -10160 240
rect -10140 220 -10070 240
rect -10050 220 -9980 240
rect -9960 220 -9890 240
rect -9870 220 -9800 240
rect -9780 220 -9710 240
rect -9690 220 -9620 240
rect -9600 220 -9530 240
rect -9510 220 -9440 240
rect -9420 220 -9350 240
rect -9330 220 -9260 240
rect -9240 220 -9170 240
rect -9150 220 -9080 240
rect -9060 220 -8990 240
rect -8970 220 -8900 240
rect -8880 220 -8810 240
rect -8790 220 -8720 240
rect -8700 220 -8630 240
rect -8610 220 -8540 240
rect -8520 220 -8450 240
rect -8430 220 -8360 240
rect -8340 220 -8270 240
rect -8250 220 -8180 240
rect -8160 220 -8090 240
rect -8070 220 -8000 240
rect -7980 220 -7910 240
rect -7890 220 -7820 240
rect -7800 220 -7730 240
rect -7710 220 -7640 240
rect -7620 220 -7550 240
rect -7530 220 -7460 240
rect -7440 220 -7370 240
rect -7350 220 -7280 240
rect -7260 220 -7190 240
rect -7170 220 -7100 240
rect -7080 220 -7010 240
rect -6990 220 -6920 240
rect -6900 220 -6830 240
rect -6810 220 -6740 240
rect -6720 220 -6650 240
rect -6630 220 -6560 240
rect -6540 220 -6470 240
rect -6450 220 -6380 240
rect -6360 220 -6290 240
rect -6270 220 -6200 240
rect -6180 220 -6110 240
rect -6090 220 -6020 240
rect -6000 220 -5930 240
rect -5910 220 -5840 240
rect -5820 220 -5750 240
rect -5730 220 -5660 240
rect -5640 220 -5570 240
rect -5550 220 -5480 240
rect -5460 220 -5390 240
rect -5370 220 -5300 240
rect -5280 220 -5210 240
rect -5190 220 -5120 240
rect -5100 220 -5030 240
rect -5010 220 -4940 240
rect -4920 220 -4850 240
rect -4830 220 -4760 240
rect -4740 220 -4670 240
rect -4650 220 -4580 240
rect -4560 220 -4490 240
rect -4470 220 -4400 240
rect -4380 220 -4310 240
rect -4290 220 -4220 240
rect -4200 220 -4130 240
rect -4110 220 -4040 240
rect -4020 220 -3950 240
rect -3930 220 -3860 240
rect -3840 220 -3770 240
rect -3750 220 -3680 240
rect -3660 220 -3590 240
rect -3570 220 -3500 240
rect -3480 220 -3410 240
rect -3390 220 -3320 240
rect -3300 220 -3230 240
rect -3210 220 -3140 240
rect -3120 220 -3050 240
rect -3030 220 -2960 240
rect -2940 220 -2870 240
rect -2850 220 -2780 240
rect -2760 220 -2690 240
rect -2670 220 -2600 240
rect -2580 220 -2510 240
rect -2490 220 -2420 240
rect -2400 220 -2330 240
rect -2310 220 -2240 240
rect -2220 220 -2150 240
rect -2130 220 -2060 240
rect -2040 220 -1970 240
rect -1950 220 -1880 240
rect -1860 220 -1790 240
rect -1770 220 -1700 240
rect -1680 220 -1610 240
rect -1590 220 -1520 240
rect -1500 220 -1430 240
rect -1410 220 -1340 240
rect -1320 220 -1250 240
rect -1230 220 -1160 240
rect -1140 220 -1070 240
rect -1050 220 -980 240
rect -960 220 -890 240
rect -870 220 -800 240
rect -780 220 -710 240
rect -690 220 -620 240
rect -600 220 -530 240
rect -510 220 -440 240
rect -420 220 -350 240
rect -330 220 -260 240
rect -240 220 -170 240
rect -150 220 -80 240
rect -60 220 120 240
rect -11690 20 -11670 220
rect -11520 175 -11510 195
rect -11490 175 -11420 195
rect -11400 175 -11330 195
rect -11310 175 -11240 195
rect -11220 175 -11150 195
rect -11130 175 -11060 195
rect -11040 175 -10970 195
rect -10950 175 -10880 195
rect -10860 175 -10850 195
rect -10800 175 -10790 195
rect -10770 175 -10700 195
rect -10680 175 -10670 195
rect -10620 175 -10610 195
rect -10590 175 -10520 195
rect -10500 175 -10490 195
rect -10440 175 -10430 195
rect -10410 175 -10340 195
rect -10320 175 -10310 195
rect -10260 175 -10250 195
rect -10230 175 -10160 195
rect -10140 175 -10130 195
rect -10080 175 -10070 195
rect -10050 175 -9980 195
rect -9960 175 -9890 195
rect -9870 175 -9800 195
rect -9780 175 -9710 195
rect -9690 175 -9620 195
rect -9600 175 -9530 195
rect -9510 175 -9440 195
rect -9420 175 -9350 195
rect -9330 175 -9260 195
rect -9240 175 -9170 195
rect -9150 175 -9080 195
rect -9060 175 -8990 195
rect -8970 175 -8900 195
rect -8880 175 -8810 195
rect -8790 175 -8720 195
rect -8700 175 -8630 195
rect -8610 175 -8540 195
rect -8520 175 -8450 195
rect -8430 175 -8360 195
rect -8340 175 -8270 195
rect -8250 175 -8180 195
rect -8160 175 -8090 195
rect -8070 175 -8000 195
rect -7980 175 -7970 195
rect -7920 175 -7910 195
rect -7890 175 -7820 195
rect -7800 175 -7790 195
rect -7740 175 -7730 195
rect -7710 175 -7640 195
rect -7620 175 -7610 195
rect -7560 175 -7550 195
rect -7530 175 -7460 195
rect -7440 175 -7430 195
rect -7380 175 -7370 195
rect -7350 175 -7280 195
rect -7260 175 -7250 195
rect -7200 175 -7190 195
rect -7170 175 -7100 195
rect -7080 175 -7070 195
rect -7020 175 -7010 195
rect -6990 175 -6920 195
rect -6900 175 -6890 195
rect -6840 175 -6830 195
rect -6810 175 -6740 195
rect -6720 175 -6710 195
rect -6660 175 -6650 195
rect -6630 175 -6560 195
rect -6540 175 -6530 195
rect -6480 175 -6470 195
rect -6450 175 -6380 195
rect -6360 175 -6290 195
rect -6270 175 -6200 195
rect -6180 175 -6110 195
rect -6090 175 -6020 195
rect -6000 175 -5930 195
rect -5910 175 -5840 195
rect -5820 175 -5750 195
rect -5730 175 -5660 195
rect -5640 175 -5570 195
rect -5550 175 -5480 195
rect -5460 175 -5390 195
rect -5370 175 -5300 195
rect -5280 175 -5210 195
rect -5190 175 -5120 195
rect -5100 175 -5030 195
rect -5010 175 -4940 195
rect -4920 175 -4850 195
rect -4830 175 -4760 195
rect -4740 175 -4670 195
rect -4650 175 -4580 195
rect -4560 175 -4490 195
rect -4470 175 -4400 195
rect -4380 175 -4370 195
rect -4320 175 -4310 195
rect -4290 175 -4220 195
rect -4200 175 -4190 195
rect -4140 175 -4130 195
rect -4110 175 -4040 195
rect -4020 175 -4010 195
rect -3960 175 -3950 195
rect -3930 175 -3860 195
rect -3840 175 -3830 195
rect -3780 175 -3770 195
rect -3750 175 -3680 195
rect -3660 175 -3650 195
rect -3600 175 -3590 195
rect -3570 175 -3500 195
rect -3480 175 -3470 195
rect -3420 175 -3410 195
rect -3390 175 -3320 195
rect -3300 175 -3290 195
rect -3240 175 -3230 195
rect -3210 175 -3140 195
rect -3120 175 -3110 195
rect -3060 175 -3050 195
rect -3030 175 -2960 195
rect -2940 175 -2930 195
rect -2880 175 -2870 195
rect -2850 175 -2780 195
rect -2760 175 -2750 195
rect -2700 175 -2690 195
rect -2670 175 -2600 195
rect -2580 175 -2570 195
rect -2520 175 -2510 195
rect -2490 175 -2420 195
rect -2400 175 -2390 195
rect -2340 175 -2330 195
rect -2310 175 -2240 195
rect -2220 175 -2210 195
rect -2160 175 -2150 195
rect -2130 175 -2060 195
rect -2040 175 -2030 195
rect -1980 175 -1970 195
rect -1950 175 -1880 195
rect -1860 175 -1850 195
rect -1800 175 -1790 195
rect -1770 175 -1700 195
rect -1680 175 -1670 195
rect -1620 175 -1610 195
rect -1590 175 -1520 195
rect -1500 175 -1490 195
rect -1440 175 -1430 195
rect -1410 175 -1340 195
rect -1320 175 -1310 195
rect -1260 175 -1250 195
rect -1230 175 -1160 195
rect -1140 175 -1130 195
rect -1080 175 -1070 195
rect -1050 175 -980 195
rect -960 175 -950 195
rect -900 175 -890 195
rect -870 175 -800 195
rect -780 175 -770 195
rect -720 175 -710 195
rect -690 175 -620 195
rect -600 175 -530 195
rect -510 175 -440 195
rect -420 175 -350 195
rect -330 175 -260 195
rect -240 175 -170 195
rect -150 175 -80 195
rect -60 175 -50 195
rect -11555 140 -11535 150
rect -11555 50 -11535 60
rect -11465 140 -11445 150
rect -11465 50 -11445 60
rect -11375 140 -11355 150
rect -11375 50 -11355 60
rect -11285 140 -11265 175
rect -11285 50 -11265 60
rect -11195 140 -11175 150
rect -11195 50 -11175 60
rect -11105 140 -11085 175
rect -11105 50 -11085 60
rect -11015 140 -10995 150
rect -11015 50 -10995 60
rect -10925 140 -10905 150
rect -10925 50 -10905 60
rect -10835 140 -10815 150
rect -10835 50 -10815 60
rect -10745 140 -10725 150
rect -10745 50 -10725 60
rect -10655 140 -10635 150
rect -10655 50 -10635 60
rect -10565 140 -10545 150
rect -10565 50 -10545 60
rect -10475 140 -10455 150
rect -10475 50 -10455 60
rect -10385 140 -10365 150
rect -10385 50 -10365 60
rect -10295 140 -10275 150
rect -10295 50 -10275 60
rect -10205 140 -10185 150
rect -10205 50 -10185 60
rect -10115 140 -10095 150
rect -10115 50 -10095 60
rect -10025 140 -10005 150
rect -10025 50 -10005 60
rect -9935 140 -9915 150
rect -9935 50 -9915 60
rect -9845 140 -9825 150
rect -9845 50 -9825 60
rect -9755 140 -9735 150
rect -9755 50 -9735 60
rect -9665 140 -9645 150
rect -9665 50 -9645 60
rect -9575 140 -9555 150
rect -9575 50 -9555 60
rect -9485 140 -9465 150
rect -9485 50 -9465 60
rect -9395 140 -9375 150
rect -9395 50 -9375 60
rect -9305 140 -9285 150
rect -9305 50 -9285 60
rect -9215 140 -9195 150
rect -9215 50 -9195 60
rect -9125 140 -9105 150
rect -9125 50 -9105 60
rect -9035 140 -9015 175
rect -9035 50 -9015 60
rect -8945 140 -8925 150
rect -8945 50 -8925 60
rect -8855 140 -8835 150
rect -8855 50 -8835 60
rect -8765 140 -8745 150
rect -8765 50 -8745 60
rect -8675 140 -8655 150
rect -8675 50 -8655 60
rect -8585 140 -8565 150
rect -8585 50 -8565 60
rect -8495 140 -8475 150
rect -8495 50 -8475 60
rect -8405 140 -8385 150
rect -8405 50 -8385 60
rect -8315 140 -8295 150
rect -8315 50 -8295 60
rect -8225 140 -8205 150
rect -8225 50 -8205 60
rect -8135 140 -8115 150
rect -8135 50 -8115 60
rect -8045 140 -8025 150
rect -8045 50 -8025 60
rect -7955 140 -7935 150
rect -7955 50 -7935 60
rect -7865 140 -7845 150
rect -7865 50 -7845 60
rect -7775 140 -7755 150
rect -7775 50 -7755 60
rect -7685 140 -7665 150
rect -7685 50 -7665 60
rect -7595 140 -7575 150
rect -7595 50 -7575 60
rect -7505 140 -7485 150
rect -7505 50 -7485 60
rect -7415 140 -7395 150
rect -7415 50 -7395 60
rect -7325 140 -7305 150
rect -7325 50 -7305 60
rect -7235 140 -7215 150
rect -7235 50 -7215 60
rect -7145 140 -7125 150
rect -7145 50 -7125 60
rect -7055 140 -7035 150
rect -7055 50 -7035 60
rect -6965 140 -6945 150
rect -6965 50 -6945 60
rect -6875 140 -6855 150
rect -6875 50 -6855 60
rect -6785 140 -6765 150
rect -6785 50 -6765 60
rect -6695 140 -6675 150
rect -6695 50 -6675 60
rect -6605 140 -6585 150
rect -6605 50 -6585 60
rect -6515 140 -6495 150
rect -6515 50 -6495 60
rect -6425 140 -6405 150
rect -6425 50 -6405 60
rect -6335 140 -6315 150
rect -6335 50 -6315 60
rect -6245 140 -6225 150
rect -6245 50 -6225 60
rect -6155 140 -6135 150
rect -6155 50 -6135 60
rect -6065 140 -6045 150
rect -6065 50 -6045 60
rect -5975 140 -5955 150
rect -5975 50 -5955 60
rect -5885 140 -5865 150
rect -5885 50 -5865 60
rect -5795 140 -5775 150
rect -5795 50 -5775 60
rect -5705 140 -5685 150
rect -5705 50 -5685 60
rect -5615 140 -5595 150
rect -5615 50 -5595 60
rect -5525 140 -5505 150
rect -5525 50 -5505 60
rect -5435 140 -5415 175
rect -5435 50 -5415 60
rect -5345 140 -5325 150
rect -5345 50 -5325 60
rect -5255 140 -5235 150
rect -5255 50 -5235 60
rect -5165 140 -5145 150
rect -5165 50 -5145 60
rect -5075 140 -5055 150
rect -5075 50 -5055 60
rect -4985 140 -4965 150
rect -4985 50 -4965 60
rect -4895 140 -4875 150
rect -4895 50 -4875 60
rect -4805 140 -4785 150
rect -4805 50 -4785 60
rect -4715 140 -4695 150
rect -4715 50 -4695 60
rect -4625 140 -4605 150
rect -4625 50 -4605 60
rect -4535 140 -4515 150
rect -4535 50 -4515 60
rect -4445 140 -4425 150
rect -4445 50 -4425 60
rect -4355 140 -4335 150
rect -4355 50 -4335 60
rect -4265 140 -4245 150
rect -4265 50 -4245 60
rect -4175 140 -4155 150
rect -4175 50 -4155 60
rect -4085 140 -4065 150
rect -4085 50 -4065 60
rect -3995 140 -3975 150
rect -3995 50 -3975 60
rect -3905 140 -3885 150
rect -3905 50 -3885 60
rect -3815 140 -3795 150
rect -3815 50 -3795 60
rect -3725 140 -3705 150
rect -3725 50 -3705 60
rect -3635 140 -3615 150
rect -3635 50 -3615 60
rect -3545 140 -3525 150
rect -3545 50 -3525 60
rect -3455 140 -3435 150
rect -3455 50 -3435 60
rect -3365 140 -3345 150
rect -3365 50 -3345 60
rect -3275 140 -3255 150
rect -3275 50 -3255 60
rect -3185 140 -3165 150
rect -3185 50 -3165 60
rect -3095 140 -3075 150
rect -3095 50 -3075 60
rect -3005 140 -2985 150
rect -3005 50 -2985 60
rect -2915 140 -2895 150
rect -2915 50 -2895 60
rect -2825 140 -2805 150
rect -2825 50 -2805 60
rect -2735 140 -2715 150
rect -2735 50 -2715 60
rect -2645 140 -2625 150
rect -2645 50 -2625 60
rect -2555 140 -2535 150
rect -2555 50 -2535 60
rect -2465 140 -2445 150
rect -2465 50 -2445 60
rect -2375 140 -2355 150
rect -2375 50 -2355 60
rect -2285 140 -2265 150
rect -2285 50 -2265 60
rect -2195 140 -2175 150
rect -2195 50 -2175 60
rect -2105 140 -2085 150
rect -2105 50 -2085 60
rect -2015 140 -1995 150
rect -2015 50 -1995 60
rect -1925 140 -1905 150
rect -1925 50 -1905 60
rect -1835 140 -1815 150
rect -1835 50 -1815 60
rect -1745 140 -1725 150
rect -1745 50 -1725 60
rect -1655 140 -1635 150
rect -1655 50 -1635 60
rect -1565 140 -1545 150
rect -1565 50 -1545 60
rect -1475 140 -1455 150
rect -1475 50 -1455 60
rect -1385 140 -1365 150
rect -1385 50 -1365 60
rect -1295 140 -1275 150
rect -1295 50 -1275 60
rect -1205 140 -1185 150
rect -1205 50 -1185 60
rect -1115 140 -1095 150
rect -1115 50 -1095 60
rect -1025 140 -1005 150
rect -1025 50 -1005 60
rect -935 140 -915 150
rect -935 50 -915 60
rect -845 140 -825 150
rect -845 50 -825 60
rect -755 140 -735 150
rect -755 50 -735 60
rect -665 140 -645 150
rect -665 50 -645 60
rect -575 140 -555 150
rect -575 50 -555 60
rect -485 140 -465 175
rect -485 50 -465 60
rect -395 140 -375 150
rect -395 50 -375 60
rect -305 140 -285 175
rect -305 50 -285 60
rect -215 140 -195 150
rect -215 50 -195 60
rect -125 140 -105 150
rect -125 50 -105 60
rect -35 140 -15 150
rect -35 50 -15 60
rect 100 20 120 220
rect -11700 0 -11690 20
rect -11670 0 -11555 20
rect -11535 0 -11510 20
rect -11490 0 -11420 20
rect -11400 0 -11330 20
rect -11310 0 -11240 20
rect -11220 0 -11150 20
rect -11130 0 -11060 20
rect -11040 0 -10970 20
rect -10950 0 -10880 20
rect -10860 0 -10835 20
rect -10815 0 -10790 20
rect -10770 0 -10700 20
rect -10680 0 -10655 20
rect -10635 0 -10610 20
rect -10590 0 -10520 20
rect -10500 0 -10475 20
rect -10455 0 -10430 20
rect -10410 0 -10340 20
rect -10320 0 -10295 20
rect -10275 0 -10250 20
rect -10230 0 -10160 20
rect -10140 0 -10115 20
rect -10095 0 -10070 20
rect -10050 0 -9980 20
rect -9960 0 -9935 20
rect -9915 0 -9890 20
rect -9870 0 -9800 20
rect -9780 0 -9755 20
rect -9735 0 -9710 20
rect -9690 0 -9620 20
rect -9600 0 -9575 20
rect -9555 0 -9530 20
rect -9510 0 -9440 20
rect -9420 0 -9395 20
rect -9375 0 -9350 20
rect -9330 0 -9260 20
rect -9240 0 -9215 20
rect -9195 0 -9170 20
rect -9150 0 -9080 20
rect -9060 0 -9035 20
rect -9015 0 -8990 20
rect -8970 0 -8900 20
rect -8880 0 -8855 20
rect -8835 0 -8810 20
rect -8790 0 -8720 20
rect -8700 0 -8675 20
rect -8655 0 -8630 20
rect -8610 0 -8540 20
rect -8520 0 -8495 20
rect -8475 0 -8450 20
rect -8430 0 -8360 20
rect -8340 0 -8315 20
rect -8295 0 -8270 20
rect -8250 0 -8180 20
rect -8160 0 -8135 20
rect -8115 0 -8090 20
rect -8070 0 -8000 20
rect -7980 0 -7955 20
rect -7935 0 -7910 20
rect -7890 0 -7820 20
rect -7800 0 -7775 20
rect -7755 0 -7730 20
rect -7710 0 -7640 20
rect -7620 0 -7595 20
rect -7575 0 -7550 20
rect -7530 0 -7460 20
rect -7440 0 -7415 20
rect -7395 0 -7370 20
rect -7350 0 -7280 20
rect -7260 0 -7235 20
rect -7215 0 -7190 20
rect -7170 0 -7100 20
rect -7080 0 -7055 20
rect -7035 0 -7010 20
rect -6990 0 -6920 20
rect -6900 0 -6875 20
rect -6855 0 -6830 20
rect -6810 0 -6740 20
rect -6720 0 -6695 20
rect -6675 0 -6650 20
rect -6630 0 -6560 20
rect -6540 0 -6515 20
rect -6495 0 -6470 20
rect -6450 0 -6380 20
rect -6360 0 -6335 20
rect -6315 0 -6290 20
rect -6270 0 -6200 20
rect -6180 0 -6155 20
rect -6135 0 -6110 20
rect -6090 0 -6020 20
rect -6000 0 -5975 20
rect -5955 0 -5930 20
rect -5910 0 -5840 20
rect -5820 0 -5795 20
rect -5775 0 -5750 20
rect -5730 0 -5660 20
rect -5640 0 -5615 20
rect -5595 0 -5570 20
rect -5550 0 -5480 20
rect -5460 0 -5435 20
rect -5415 0 -5390 20
rect -5370 0 -5300 20
rect -5280 0 -5255 20
rect -5235 0 -5210 20
rect -5190 0 -5120 20
rect -5100 0 -5075 20
rect -5055 0 -5030 20
rect -5010 0 -4940 20
rect -4920 0 -4895 20
rect -4875 0 -4850 20
rect -4830 0 -4760 20
rect -4740 0 -4715 20
rect -4695 0 -4670 20
rect -4650 0 -4580 20
rect -4560 0 -4535 20
rect -4515 0 -4490 20
rect -4470 0 -4400 20
rect -4380 0 -4355 20
rect -4335 0 -4310 20
rect -4290 0 -4220 20
rect -4200 0 -4175 20
rect -4155 0 -4130 20
rect -4110 0 -4040 20
rect -4020 0 -3995 20
rect -3975 0 -3950 20
rect -3930 0 -3860 20
rect -3840 0 -3815 20
rect -3795 0 -3770 20
rect -3750 0 -3680 20
rect -3660 0 -3635 20
rect -3615 0 -3590 20
rect -3570 0 -3500 20
rect -3480 0 -3455 20
rect -3435 0 -3410 20
rect -3390 0 -3320 20
rect -3300 0 -3275 20
rect -3255 0 -3230 20
rect -3210 0 -3140 20
rect -3120 0 -3095 20
rect -3075 0 -3050 20
rect -3030 0 -2960 20
rect -2940 0 -2915 20
rect -2895 0 -2870 20
rect -2850 0 -2780 20
rect -2760 0 -2735 20
rect -2715 0 -2690 20
rect -2670 0 -2600 20
rect -2580 0 -2555 20
rect -2535 0 -2510 20
rect -2490 0 -2420 20
rect -2400 0 -2375 20
rect -2355 0 -2330 20
rect -2310 0 -2240 20
rect -2220 0 -2195 20
rect -2175 0 -2150 20
rect -2130 0 -2060 20
rect -2040 0 -2015 20
rect -1995 0 -1970 20
rect -1950 0 -1880 20
rect -1860 0 -1835 20
rect -1815 0 -1790 20
rect -1770 0 -1700 20
rect -1680 0 -1655 20
rect -1635 0 -1610 20
rect -1590 0 -1520 20
rect -1500 0 -1475 20
rect -1455 0 -1430 20
rect -1410 0 -1340 20
rect -1320 0 -1295 20
rect -1275 0 -1250 20
rect -1230 0 -1160 20
rect -1140 0 -1115 20
rect -1095 0 -1070 20
rect -1050 0 -980 20
rect -960 0 -935 20
rect -915 0 -890 20
rect -870 0 -800 20
rect -780 0 -755 20
rect -735 0 -710 20
rect -690 0 -620 20
rect -600 0 -530 20
rect -510 0 -440 20
rect -420 0 -350 20
rect -330 0 -260 20
rect -240 0 -170 20
rect -150 0 -80 20
rect -60 0 -35 20
rect -15 0 100 20
rect 120 0 130 20
<< viali >>
rect -11690 1975 -11670 1995
rect -11555 1975 -11535 1995
rect -10835 1975 -10815 1995
rect -10655 1975 -10635 1995
rect -10475 1975 -10455 1995
rect -10295 1975 -10275 1995
rect -10115 1975 -10095 1995
rect -9935 1975 -9915 1995
rect -9755 1975 -9735 1995
rect -9575 1975 -9555 1995
rect -9395 1975 -9375 1995
rect -9215 1975 -9195 1995
rect -9035 1975 -9015 1995
rect -8855 1975 -8835 1995
rect -8675 1975 -8655 1995
rect -8495 1975 -8475 1995
rect -8315 1975 -8295 1995
rect -8135 1975 -8115 1995
rect -7955 1975 -7935 1995
rect -7775 1975 -7755 1995
rect -7595 1975 -7575 1995
rect -7415 1975 -7395 1995
rect -7235 1975 -7215 1995
rect -7055 1975 -7035 1995
rect -6875 1975 -6855 1995
rect -6695 1975 -6675 1995
rect -6515 1975 -6495 1995
rect -6335 1975 -6315 1995
rect -6155 1975 -6135 1995
rect -5975 1975 -5955 1995
rect -5795 1975 -5775 1995
rect -5615 1975 -5595 1995
rect -5435 1975 -5415 1995
rect -5255 1975 -5235 1995
rect -5075 1975 -5055 1995
rect -4895 1975 -4875 1995
rect -4715 1975 -4695 1995
rect -4535 1975 -4515 1995
rect -4355 1975 -4335 1995
rect -4175 1975 -4155 1995
rect -3995 1975 -3975 1995
rect -3815 1975 -3795 1995
rect -3635 1975 -3615 1995
rect -3455 1975 -3435 1995
rect -3275 1975 -3255 1995
rect -3095 1975 -3075 1995
rect -2915 1975 -2895 1995
rect -2735 1975 -2715 1995
rect -2555 1975 -2535 1995
rect -2375 1975 -2355 1995
rect -2195 1975 -2175 1995
rect -2015 1975 -1995 1995
rect -1835 1975 -1815 1995
rect -1655 1975 -1635 1995
rect -1475 1975 -1455 1995
rect -1295 1975 -1275 1995
rect -1115 1975 -1095 1995
rect -935 1975 -915 1995
rect -755 1975 -735 1995
rect -35 1975 -15 1995
rect 100 1975 120 1995
rect -11555 1855 -11535 1935
rect -10835 1855 -10815 1935
rect -10745 1855 -10725 1935
rect -10655 1855 -10635 1935
rect -10565 1855 -10545 1935
rect -10475 1855 -10455 1935
rect -10385 1855 -10365 1935
rect -10295 1855 -10275 1935
rect -10205 1855 -10185 1935
rect -10115 1855 -10095 1935
rect -10025 1855 -10005 1935
rect -9935 1855 -9915 1935
rect -9845 1855 -9825 1935
rect -9755 1855 -9735 1935
rect -9665 1855 -9645 1935
rect -9575 1855 -9555 1935
rect -9485 1855 -9465 1935
rect -9395 1855 -9375 1935
rect -9305 1855 -9285 1935
rect -9215 1855 -9195 1935
rect -9125 1855 -9105 1935
rect -9035 1855 -9015 1935
rect -8945 1855 -8925 1935
rect -8855 1855 -8835 1935
rect -8765 1855 -8745 1935
rect -8675 1855 -8655 1935
rect -8585 1855 -8565 1935
rect -8495 1855 -8475 1935
rect -8405 1855 -8385 1935
rect -8315 1855 -8295 1935
rect -8225 1855 -8205 1935
rect -8135 1855 -8115 1935
rect -8045 1855 -8025 1935
rect -7955 1855 -7935 1935
rect -7865 1855 -7845 1935
rect -7775 1855 -7755 1935
rect -7685 1855 -7665 1935
rect -7595 1855 -7575 1935
rect -7505 1855 -7485 1935
rect -7415 1855 -7395 1935
rect -7325 1855 -7305 1935
rect -7235 1855 -7215 1935
rect -7145 1855 -7125 1935
rect -7055 1855 -7035 1935
rect -6965 1855 -6945 1935
rect -6875 1855 -6855 1935
rect -6785 1855 -6765 1935
rect -6695 1855 -6675 1935
rect -6605 1855 -6585 1935
rect -6515 1855 -6495 1935
rect -6425 1855 -6405 1935
rect -6335 1855 -6315 1935
rect -6245 1855 -6225 1935
rect -6155 1855 -6135 1935
rect -6065 1855 -6045 1935
rect -5975 1855 -5955 1935
rect -5885 1855 -5865 1935
rect -5795 1855 -5775 1935
rect -5705 1855 -5685 1935
rect -5615 1855 -5595 1935
rect -5525 1855 -5505 1935
rect -5435 1855 -5415 1935
rect -5345 1855 -5325 1935
rect -5255 1855 -5235 1935
rect -5165 1855 -5145 1935
rect -5075 1855 -5055 1935
rect -4985 1855 -4965 1935
rect -4895 1855 -4875 1935
rect -4805 1855 -4785 1935
rect -4715 1855 -4695 1935
rect -4625 1855 -4605 1935
rect -4535 1855 -4515 1935
rect -4445 1855 -4425 1935
rect -4355 1855 -4335 1935
rect -4265 1855 -4245 1935
rect -4175 1855 -4155 1935
rect -4085 1855 -4065 1935
rect -3995 1855 -3975 1935
rect -3905 1855 -3885 1935
rect -3815 1855 -3795 1935
rect -3725 1855 -3705 1935
rect -3635 1855 -3615 1935
rect -3545 1855 -3525 1935
rect -3455 1855 -3435 1935
rect -3365 1855 -3345 1935
rect -3275 1855 -3255 1935
rect -3185 1855 -3165 1935
rect -3095 1855 -3075 1935
rect -3005 1855 -2985 1935
rect -2915 1855 -2895 1935
rect -2825 1855 -2805 1935
rect -2735 1855 -2715 1935
rect -2645 1855 -2625 1935
rect -2555 1855 -2535 1935
rect -2465 1855 -2445 1935
rect -2375 1855 -2355 1935
rect -2285 1855 -2265 1935
rect -2195 1855 -2175 1935
rect -2105 1855 -2085 1935
rect -2015 1855 -1995 1935
rect -1925 1855 -1905 1935
rect -1835 1855 -1815 1935
rect -1745 1855 -1725 1935
rect -1655 1855 -1635 1935
rect -1565 1855 -1545 1935
rect -1475 1855 -1455 1935
rect -1385 1855 -1365 1935
rect -1295 1855 -1275 1935
rect -1205 1855 -1185 1935
rect -1115 1855 -1095 1935
rect -1025 1855 -1005 1935
rect -935 1855 -915 1935
rect -845 1855 -825 1935
rect -755 1855 -735 1935
rect -35 1855 -15 1935
rect -10700 1800 -10680 1820
rect -10520 1800 -10500 1820
rect -10340 1800 -10320 1820
rect -10160 1800 -10140 1820
rect -9980 1800 -9960 1820
rect -9800 1800 -9780 1820
rect -9620 1800 -9600 1820
rect -9440 1800 -9420 1820
rect -9260 1800 -9240 1820
rect -9080 1800 -9060 1820
rect -8900 1800 -8880 1820
rect -8720 1800 -8700 1820
rect -8540 1800 -8520 1820
rect -8360 1800 -8340 1820
rect -8180 1800 -8160 1820
rect -8000 1800 -7980 1820
rect -7820 1800 -7800 1820
rect -7640 1800 -7620 1820
rect -7460 1800 -7440 1820
rect -7280 1800 -7260 1820
rect -7100 1800 -7080 1820
rect -6920 1800 -6900 1820
rect -6740 1800 -6720 1820
rect -6560 1800 -6540 1820
rect -6380 1800 -6360 1820
rect -6200 1800 -6180 1820
rect -6020 1800 -6000 1820
rect -5840 1800 -5820 1820
rect -5660 1800 -5640 1820
rect -5480 1800 -5460 1820
rect -5300 1800 -5280 1820
rect -5120 1800 -5100 1820
rect -4940 1800 -4920 1820
rect -4760 1800 -4740 1820
rect -4580 1800 -4560 1820
rect -4400 1800 -4380 1820
rect -4220 1800 -4200 1820
rect -4040 1800 -4020 1820
rect -3860 1800 -3840 1820
rect -3680 1800 -3660 1820
rect -3500 1800 -3480 1820
rect -3320 1800 -3300 1820
rect -3140 1800 -3120 1820
rect -2960 1800 -2940 1820
rect -2780 1800 -2760 1820
rect -2600 1800 -2580 1820
rect -2420 1800 -2400 1820
rect -2240 1800 -2220 1820
rect -2060 1800 -2040 1820
rect -1880 1800 -1860 1820
rect -1700 1800 -1680 1820
rect -1520 1800 -1500 1820
rect -1340 1800 -1320 1820
rect -1160 1800 -1140 1820
rect -980 1800 -960 1820
rect -800 1800 -780 1820
rect -10700 1715 -10680 1735
rect -10520 1715 -10500 1735
rect -9620 1715 -9600 1735
rect -9440 1715 -9420 1735
rect -9260 1715 -9240 1735
rect -9080 1715 -9060 1735
rect -8180 1715 -8160 1735
rect -8000 1715 -7980 1735
rect -7820 1715 -7800 1735
rect -7640 1715 -7620 1735
rect -4580 1715 -4560 1735
rect -4400 1715 -4380 1735
rect -4220 1715 -4200 1735
rect -4040 1715 -4020 1735
rect -980 1715 -960 1735
rect -800 1715 -780 1735
rect -125 1715 -105 1735
rect -10340 1675 -10320 1695
rect -10160 1675 -10140 1695
rect -9980 1675 -9960 1695
rect -9800 1675 -9780 1695
rect -8900 1675 -8880 1695
rect -8720 1675 -8700 1695
rect -8540 1675 -8520 1695
rect -8360 1675 -8340 1695
rect -7460 1675 -7440 1695
rect -7280 1675 -7260 1695
rect -4940 1675 -4920 1695
rect -4760 1675 -4740 1695
rect -3860 1675 -3840 1695
rect -3680 1675 -3660 1695
rect -1340 1675 -1320 1695
rect -1160 1675 -1140 1695
rect -215 1675 -195 1695
rect -11105 1635 -11085 1655
rect -9035 1635 -9015 1655
rect -8315 1635 -8295 1655
rect -3995 1635 -3975 1655
rect -3545 1635 -3525 1655
rect -3365 1635 -3345 1655
rect -3185 1635 -3165 1655
rect -3005 1635 -2985 1655
rect -2825 1635 -2805 1655
rect -2645 1635 -2625 1655
rect -2465 1635 -2445 1655
rect -2285 1635 -2265 1655
rect -2105 1635 -2085 1655
rect -1925 1635 -1905 1655
rect -1745 1635 -1725 1655
rect -1565 1635 -1545 1655
rect -1115 1635 -1095 1655
rect -11195 1595 -11175 1615
rect -10475 1595 -10455 1615
rect -9755 1595 -9735 1615
rect -7595 1595 -7575 1615
rect -7145 1595 -7125 1615
rect -6965 1595 -6945 1615
rect -6785 1595 -6765 1615
rect -6605 1595 -6585 1615
rect -6425 1595 -6405 1615
rect -6245 1595 -6225 1615
rect -6065 1595 -6045 1615
rect -5885 1595 -5865 1615
rect -5705 1595 -5685 1615
rect -5525 1595 -5505 1615
rect -5345 1595 -5325 1615
rect -5165 1595 -5145 1615
rect -4715 1595 -4695 1615
rect -11285 1555 -11265 1575
rect -3590 1555 -3570 1575
rect -3410 1555 -3390 1575
rect -3230 1555 -3210 1575
rect -3050 1555 -3030 1575
rect -2870 1555 -2850 1575
rect -2690 1555 -2670 1575
rect -2510 1555 -2490 1575
rect -2330 1555 -2310 1575
rect -2150 1555 -2130 1575
rect -1970 1555 -1950 1575
rect -1790 1555 -1770 1575
rect -1610 1555 -1590 1575
rect -11375 1515 -11355 1535
rect -7190 1515 -7170 1535
rect -7010 1515 -6990 1535
rect -6830 1515 -6810 1535
rect -6650 1515 -6630 1535
rect -6470 1515 -6450 1535
rect -6290 1515 -6270 1535
rect -6110 1515 -6090 1535
rect -5930 1515 -5910 1535
rect -5750 1515 -5730 1535
rect -5570 1515 -5550 1535
rect -5390 1515 -5370 1535
rect -5210 1515 -5190 1535
rect -11465 1475 -11445 1495
rect -10115 1475 -10095 1495
rect -7235 1475 -7215 1495
rect -5075 1475 -5055 1495
rect -10790 1435 -10770 1455
rect -10610 1435 -10590 1455
rect -9710 1435 -9690 1455
rect -9530 1435 -9510 1455
rect -9350 1435 -9330 1455
rect -9170 1435 -9150 1455
rect -8675 1435 -8655 1455
rect -8270 1435 -8250 1455
rect -8090 1435 -8070 1455
rect -3635 1435 -3615 1455
rect -1475 1435 -1455 1455
rect -485 1435 -465 1455
rect -10430 1395 -10410 1415
rect -10250 1395 -10230 1415
rect -10070 1395 -10050 1415
rect -9890 1395 -9870 1415
rect -8990 1395 -8970 1415
rect -8810 1395 -8790 1415
rect -8630 1395 -8610 1415
rect -8450 1395 -8430 1415
rect -7550 1395 -7530 1415
rect -7370 1395 -7350 1415
rect -5030 1395 -5010 1415
rect -4850 1395 -4830 1415
rect -3950 1395 -3930 1415
rect -3770 1395 -3750 1415
rect -1430 1395 -1410 1415
rect -1250 1395 -1230 1415
rect -305 1395 -285 1415
rect -7910 1355 -7890 1375
rect -7730 1355 -7710 1375
rect -4670 1355 -4650 1375
rect -4490 1355 -4470 1375
rect -4310 1355 -4290 1375
rect -4130 1355 -4110 1375
rect -1070 1355 -1050 1375
rect -890 1355 -870 1375
rect -395 1355 -375 1375
rect -7235 1275 -7215 1295
rect -7055 1275 -7035 1295
rect -6875 1275 -6855 1295
rect -6695 1275 -6675 1295
rect -6515 1275 -6495 1295
rect -6335 1275 -6315 1295
rect -6155 1275 -6135 1295
rect -5975 1275 -5955 1295
rect -5795 1275 -5775 1295
rect -5615 1275 -5595 1295
rect -5435 1275 -5415 1295
rect -5255 1275 -5235 1295
rect -5075 1275 -5055 1295
rect -3635 1275 -3615 1295
rect -3455 1275 -3435 1295
rect -3275 1275 -3255 1295
rect -3095 1275 -3075 1295
rect -2915 1275 -2895 1295
rect -2735 1275 -2715 1295
rect -2555 1275 -2535 1295
rect -2375 1275 -2355 1295
rect -2195 1275 -2175 1295
rect -2015 1275 -1995 1295
rect -1835 1275 -1815 1295
rect -1655 1275 -1635 1295
rect -1475 1275 -1455 1295
rect -575 1275 -555 1295
rect -10790 1190 -10770 1210
rect -10610 1190 -10590 1210
rect -10430 1190 -10410 1210
rect -10250 1190 -10230 1210
rect -10070 1190 -10050 1210
rect -9890 1190 -9870 1210
rect -9710 1190 -9690 1210
rect -9530 1190 -9510 1210
rect -9350 1190 -9330 1210
rect -9170 1190 -9150 1210
rect -8990 1190 -8970 1210
rect -8810 1190 -8790 1210
rect -8630 1190 -8610 1210
rect -8450 1190 -8430 1210
rect -8270 1190 -8250 1210
rect -8090 1190 -8070 1210
rect -7910 1190 -7890 1210
rect -7730 1190 -7710 1210
rect -7550 1190 -7530 1210
rect -7370 1190 -7350 1210
rect -7190 1190 -7170 1210
rect -7010 1190 -6990 1210
rect -6830 1190 -6810 1210
rect -6650 1190 -6630 1210
rect -6470 1190 -6450 1210
rect -6290 1190 -6270 1210
rect -6110 1190 -6090 1210
rect -5930 1190 -5910 1210
rect -5750 1190 -5730 1210
rect -5570 1190 -5550 1210
rect -5390 1190 -5370 1210
rect -5210 1190 -5190 1210
rect -5030 1190 -5010 1210
rect -4850 1190 -4830 1210
rect -4670 1190 -4650 1210
rect -4490 1190 -4470 1210
rect -4310 1190 -4290 1210
rect -4130 1190 -4110 1210
rect -3950 1190 -3930 1210
rect -3770 1190 -3750 1210
rect -3590 1190 -3570 1210
rect -3410 1190 -3390 1210
rect -3230 1190 -3210 1210
rect -3050 1190 -3030 1210
rect -2870 1190 -2850 1210
rect -2690 1190 -2670 1210
rect -2510 1190 -2490 1210
rect -2330 1190 -2310 1210
rect -2150 1190 -2130 1210
rect -1970 1190 -1950 1210
rect -1790 1190 -1770 1210
rect -1610 1190 -1590 1210
rect -1430 1190 -1410 1210
rect -1250 1190 -1230 1210
rect -1070 1190 -1050 1210
rect -890 1190 -870 1210
rect -11555 1075 -11535 1155
rect -10835 1075 -10815 1155
rect -10745 1075 -10725 1155
rect -10655 1075 -10635 1155
rect -10565 1075 -10545 1155
rect -10475 1075 -10455 1155
rect -10385 1075 -10365 1155
rect -10295 1075 -10275 1155
rect -10205 1075 -10185 1155
rect -10115 1075 -10095 1155
rect -10025 1075 -10005 1155
rect -9935 1075 -9915 1155
rect -9845 1075 -9825 1155
rect -9755 1075 -9735 1155
rect -9665 1075 -9645 1155
rect -9575 1075 -9555 1155
rect -9485 1075 -9465 1155
rect -9395 1075 -9375 1155
rect -9305 1075 -9285 1155
rect -9215 1075 -9195 1155
rect -9125 1075 -9105 1155
rect -9035 1075 -9015 1155
rect -8945 1075 -8925 1155
rect -8855 1075 -8835 1155
rect -8765 1075 -8745 1155
rect -8675 1075 -8655 1155
rect -8585 1075 -8565 1155
rect -8495 1075 -8475 1155
rect -8405 1075 -8385 1155
rect -8315 1075 -8295 1155
rect -8225 1075 -8205 1155
rect -8135 1075 -8115 1155
rect -8045 1075 -8025 1155
rect -7955 1075 -7935 1155
rect -7865 1075 -7845 1155
rect -7775 1075 -7755 1155
rect -7685 1075 -7665 1155
rect -7595 1075 -7575 1155
rect -7505 1075 -7485 1155
rect -7415 1075 -7395 1155
rect -7325 1075 -7305 1155
rect -7235 1075 -7215 1155
rect -7145 1075 -7125 1155
rect -7055 1075 -7035 1155
rect -6965 1075 -6945 1155
rect -6875 1075 -6855 1155
rect -6785 1075 -6765 1155
rect -6695 1075 -6675 1155
rect -6605 1075 -6585 1155
rect -6515 1075 -6495 1155
rect -6425 1075 -6405 1155
rect -6335 1075 -6315 1155
rect -6245 1075 -6225 1155
rect -6155 1075 -6135 1155
rect -6065 1075 -6045 1155
rect -5975 1075 -5955 1155
rect -5885 1075 -5865 1155
rect -5795 1075 -5775 1155
rect -5705 1075 -5685 1155
rect -5615 1075 -5595 1155
rect -5525 1075 -5505 1155
rect -5435 1075 -5415 1155
rect -5345 1075 -5325 1155
rect -5255 1075 -5235 1155
rect -5165 1075 -5145 1155
rect -5075 1075 -5055 1155
rect -4985 1075 -4965 1155
rect -4895 1075 -4875 1155
rect -4805 1075 -4785 1155
rect -4715 1075 -4695 1155
rect -4625 1075 -4605 1155
rect -4535 1075 -4515 1155
rect -4445 1075 -4425 1155
rect -4355 1075 -4335 1155
rect -4265 1075 -4245 1155
rect -4175 1075 -4155 1155
rect -4085 1075 -4065 1155
rect -3995 1075 -3975 1155
rect -3905 1075 -3885 1155
rect -3815 1075 -3795 1155
rect -3725 1075 -3705 1155
rect -3635 1075 -3615 1155
rect -3545 1075 -3525 1155
rect -3455 1075 -3435 1155
rect -3365 1075 -3345 1155
rect -3275 1075 -3255 1155
rect -3185 1075 -3165 1155
rect -3095 1075 -3075 1155
rect -3005 1075 -2985 1155
rect -2915 1075 -2895 1155
rect -2825 1075 -2805 1155
rect -2735 1075 -2715 1155
rect -2645 1075 -2625 1155
rect -2555 1075 -2535 1155
rect -2465 1075 -2445 1155
rect -2375 1075 -2355 1155
rect -2285 1075 -2265 1155
rect -2195 1075 -2175 1155
rect -2105 1075 -2085 1155
rect -2015 1075 -1995 1155
rect -1925 1075 -1905 1155
rect -1835 1075 -1815 1155
rect -1745 1075 -1725 1155
rect -1655 1075 -1635 1155
rect -1565 1075 -1545 1155
rect -1475 1075 -1455 1155
rect -1385 1075 -1365 1155
rect -1295 1075 -1275 1155
rect -1205 1075 -1185 1155
rect -1115 1075 -1095 1155
rect -1025 1075 -1005 1155
rect -935 1075 -915 1155
rect -845 1075 -825 1155
rect -755 1075 -735 1155
rect -35 1075 -15 1155
rect -11555 1015 -11535 1035
rect -10835 1015 -10815 1035
rect -10655 1015 -10635 1035
rect -10475 1015 -10455 1035
rect -10295 1015 -10275 1035
rect -10115 1015 -10095 1035
rect -9935 1015 -9915 1035
rect -9755 1015 -9735 1035
rect -9575 1015 -9555 1035
rect -9395 1015 -9375 1035
rect -9215 1015 -9195 1035
rect -9035 1015 -9015 1035
rect -8855 1015 -8835 1035
rect -8675 1015 -8655 1035
rect -8495 1015 -8475 1035
rect -8315 1015 -8295 1035
rect -8135 1015 -8115 1035
rect -7955 1015 -7935 1035
rect -7775 1015 -7755 1035
rect -7595 1015 -7575 1035
rect -7415 1015 -7395 1035
rect -7235 1015 -7215 1035
rect -7055 1015 -7035 1035
rect -6875 1015 -6855 1035
rect -6695 1015 -6675 1035
rect -6515 1015 -6495 1035
rect -6335 1015 -6315 1035
rect -6155 1015 -6135 1035
rect -5975 1015 -5955 1035
rect -5795 1015 -5775 1035
rect -5615 1015 -5595 1035
rect -5435 1015 -5415 1035
rect -5255 1015 -5235 1035
rect -5075 1015 -5055 1035
rect -4895 1015 -4875 1035
rect -4715 1015 -4695 1035
rect -4535 1015 -4515 1035
rect -4355 1015 -4335 1035
rect -4175 1015 -4155 1035
rect -3995 1015 -3975 1035
rect -3815 1015 -3795 1035
rect -3635 1015 -3615 1035
rect -3455 1015 -3435 1035
rect -3275 1015 -3255 1035
rect -3095 1015 -3075 1035
rect -2915 1015 -2895 1035
rect -2735 1015 -2715 1035
rect -2555 1015 -2535 1035
rect -2375 1015 -2355 1035
rect -2195 1015 -2175 1035
rect -2015 1015 -1995 1035
rect -1835 1015 -1815 1035
rect -1655 1015 -1635 1035
rect -1475 1015 -1455 1035
rect -1295 1015 -1275 1035
rect -1115 1015 -1095 1035
rect -935 1015 -915 1035
rect -755 1015 -735 1035
rect -35 1015 -15 1035
rect -11555 960 -11535 980
rect -10835 960 -10815 980
rect -10655 960 -10635 980
rect -10475 960 -10455 980
rect -10295 960 -10275 980
rect -10115 960 -10095 980
rect -9935 960 -9915 980
rect -9755 960 -9735 980
rect -9575 960 -9555 980
rect -9395 960 -9375 980
rect -9215 960 -9195 980
rect -9035 960 -9015 980
rect -8855 960 -8835 980
rect -8675 960 -8655 980
rect -8495 960 -8475 980
rect -8315 960 -8295 980
rect -8135 960 -8115 980
rect -7955 960 -7935 980
rect -7775 960 -7755 980
rect -7595 960 -7575 980
rect -7415 960 -7395 980
rect -7235 960 -7215 980
rect -7055 960 -7035 980
rect -6875 960 -6855 980
rect -6695 960 -6675 980
rect -6515 960 -6495 980
rect -6335 960 -6315 980
rect -6155 960 -6135 980
rect -5975 960 -5955 980
rect -5795 960 -5775 980
rect -5615 960 -5595 980
rect -5435 960 -5415 980
rect -5255 960 -5235 980
rect -5075 960 -5055 980
rect -4895 960 -4875 980
rect -4715 960 -4695 980
rect -4535 960 -4515 980
rect -4355 960 -4335 980
rect -4175 960 -4155 980
rect -3995 960 -3975 980
rect -3815 960 -3795 980
rect -3635 960 -3615 980
rect -3455 960 -3435 980
rect -3275 960 -3255 980
rect -3095 960 -3075 980
rect -2915 960 -2895 980
rect -2735 960 -2715 980
rect -2555 960 -2535 980
rect -2375 960 -2355 980
rect -2195 960 -2175 980
rect -2015 960 -1995 980
rect -1835 960 -1815 980
rect -1655 960 -1635 980
rect -1475 960 -1455 980
rect -1295 960 -1275 980
rect -1115 960 -1095 980
rect -935 960 -915 980
rect -755 960 -735 980
rect -35 960 -15 980
rect -11555 840 -11535 920
rect -10835 840 -10815 920
rect -10745 840 -10725 920
rect -10655 840 -10635 920
rect -10565 840 -10545 920
rect -10475 840 -10455 920
rect -10385 840 -10365 920
rect -10295 840 -10275 920
rect -10205 840 -10185 920
rect -10115 840 -10095 920
rect -10025 840 -10005 920
rect -9935 840 -9915 920
rect -9845 840 -9825 920
rect -9755 840 -9735 920
rect -9665 840 -9645 920
rect -9575 840 -9555 920
rect -9485 840 -9465 920
rect -9395 840 -9375 920
rect -9305 840 -9285 920
rect -9215 840 -9195 920
rect -9125 840 -9105 920
rect -9035 840 -9015 920
rect -8945 840 -8925 920
rect -8855 840 -8835 920
rect -8765 840 -8745 920
rect -8675 840 -8655 920
rect -8585 840 -8565 920
rect -8495 840 -8475 920
rect -8405 840 -8385 920
rect -8315 840 -8295 920
rect -8225 840 -8205 920
rect -8135 840 -8115 920
rect -8045 840 -8025 920
rect -7955 840 -7935 920
rect -7865 840 -7845 920
rect -7775 840 -7755 920
rect -7685 840 -7665 920
rect -7595 840 -7575 920
rect -7505 840 -7485 920
rect -7415 840 -7395 920
rect -7325 840 -7305 920
rect -7235 840 -7215 920
rect -7145 840 -7125 920
rect -7055 840 -7035 920
rect -6965 840 -6945 920
rect -6875 840 -6855 920
rect -6785 840 -6765 920
rect -6695 840 -6675 920
rect -6605 840 -6585 920
rect -6515 840 -6495 920
rect -6425 840 -6405 920
rect -6335 840 -6315 920
rect -6245 840 -6225 920
rect -6155 840 -6135 920
rect -6065 840 -6045 920
rect -5975 840 -5955 920
rect -5885 840 -5865 920
rect -5795 840 -5775 920
rect -5705 840 -5685 920
rect -5615 840 -5595 920
rect -5525 840 -5505 920
rect -5435 840 -5415 920
rect -5345 840 -5325 920
rect -5255 840 -5235 920
rect -5165 840 -5145 920
rect -5075 840 -5055 920
rect -4985 840 -4965 920
rect -4895 840 -4875 920
rect -4805 840 -4785 920
rect -4715 840 -4695 920
rect -4625 840 -4605 920
rect -4535 840 -4515 920
rect -4445 840 -4425 920
rect -4355 840 -4335 920
rect -4265 840 -4245 920
rect -4175 840 -4155 920
rect -4085 840 -4065 920
rect -3995 840 -3975 920
rect -3905 840 -3885 920
rect -3815 840 -3795 920
rect -3725 840 -3705 920
rect -3635 840 -3615 920
rect -3545 840 -3525 920
rect -3455 840 -3435 920
rect -3365 840 -3345 920
rect -3275 840 -3255 920
rect -3185 840 -3165 920
rect -3095 840 -3075 920
rect -3005 840 -2985 920
rect -2915 840 -2895 920
rect -2825 840 -2805 920
rect -2735 840 -2715 920
rect -2645 840 -2625 920
rect -2555 840 -2535 920
rect -2465 840 -2445 920
rect -2375 840 -2355 920
rect -2285 840 -2265 920
rect -2195 840 -2175 920
rect -2105 840 -2085 920
rect -2015 840 -1995 920
rect -1925 840 -1905 920
rect -1835 840 -1815 920
rect -1745 840 -1725 920
rect -1655 840 -1635 920
rect -1565 840 -1545 920
rect -1475 840 -1455 920
rect -1385 840 -1365 920
rect -1295 840 -1275 920
rect -1205 840 -1185 920
rect -1115 840 -1095 920
rect -1025 840 -1005 920
rect -935 840 -915 920
rect -845 840 -825 920
rect -755 840 -735 920
rect -35 840 -15 920
rect -10700 785 -10680 805
rect -10520 785 -10500 805
rect -10340 785 -10320 805
rect -10160 785 -10140 805
rect -9980 785 -9960 805
rect -9800 785 -9780 805
rect -9620 785 -9600 805
rect -9440 785 -9420 805
rect -9260 785 -9240 805
rect -9080 785 -9060 805
rect -8900 785 -8880 805
rect -8720 785 -8700 805
rect -8540 785 -8520 805
rect -8360 785 -8340 805
rect -8180 785 -8160 805
rect -8000 785 -7980 805
rect -7820 785 -7800 805
rect -7640 785 -7620 805
rect -7460 785 -7440 805
rect -7280 785 -7260 805
rect -7100 785 -7080 805
rect -6920 785 -6900 805
rect -6740 785 -6720 805
rect -6560 785 -6540 805
rect -6380 785 -6360 805
rect -6200 785 -6180 805
rect -6020 785 -6000 805
rect -5840 785 -5820 805
rect -5660 785 -5640 805
rect -5480 785 -5460 805
rect -5300 785 -5280 805
rect -5120 785 -5100 805
rect -4940 785 -4920 805
rect -4760 785 -4740 805
rect -4580 785 -4560 805
rect -4400 785 -4380 805
rect -4220 785 -4200 805
rect -4040 785 -4020 805
rect -3860 785 -3840 805
rect -3680 785 -3660 805
rect -3500 785 -3480 805
rect -3320 785 -3300 805
rect -3140 785 -3120 805
rect -2960 785 -2940 805
rect -2780 785 -2760 805
rect -2600 785 -2580 805
rect -2420 785 -2400 805
rect -2240 785 -2220 805
rect -2060 785 -2040 805
rect -1880 785 -1860 805
rect -1700 785 -1680 805
rect -1520 785 -1500 805
rect -1340 785 -1320 805
rect -1160 785 -1140 805
rect -980 785 -960 805
rect -800 785 -780 805
rect -10115 700 -10095 720
rect -9935 700 -9915 720
rect -9755 700 -9735 720
rect -9575 700 -9555 720
rect -9395 700 -9375 720
rect -9215 700 -9195 720
rect -9035 700 -9015 720
rect -8855 700 -8835 720
rect -8675 700 -8655 720
rect -8495 700 -8475 720
rect -8315 700 -8295 720
rect -8135 700 -8115 720
rect -7955 700 -7935 720
rect -6515 700 -6495 720
rect -6335 700 -6315 720
rect -6155 700 -6135 720
rect -5975 700 -5955 720
rect -5795 700 -5775 720
rect -5615 700 -5595 720
rect -5435 700 -5415 720
rect -5255 700 -5235 720
rect -5075 700 -5055 720
rect -4895 700 -4875 720
rect -4715 700 -4695 720
rect -4535 700 -4515 720
rect -4355 700 -4335 720
rect -575 700 -555 720
rect -10700 620 -10680 640
rect -10520 620 -10500 640
rect -7460 620 -7440 640
rect -7280 620 -7260 640
rect -7100 620 -7080 640
rect -6920 620 -6900 640
rect -3860 620 -3840 640
rect -3680 620 -3660 640
rect -395 620 -375 640
rect -10340 580 -10320 600
rect -10160 580 -10140 600
rect -7820 580 -7800 600
rect -7640 580 -7620 600
rect -6740 580 -6720 600
rect -6560 580 -6540 600
rect -4220 580 -4200 600
rect -4040 580 -4020 600
rect -3140 580 -3120 600
rect -2960 580 -2940 600
rect -2780 580 -2760 600
rect -2600 580 -2580 600
rect -1700 580 -1680 600
rect -1520 580 -1500 600
rect -1340 580 -1320 600
rect -1160 580 -1140 600
rect -305 580 -285 600
rect -10115 540 -10095 560
rect -7955 540 -7935 560
rect -3500 540 -3480 560
rect -3320 540 -3300 560
rect -2915 540 -2895 560
rect -2420 540 -2400 560
rect -2240 540 -2220 560
rect -2060 540 -2040 560
rect -1880 540 -1860 560
rect -980 540 -960 560
rect -800 540 -780 560
rect -485 540 -465 560
rect -11465 500 -11445 520
rect -6515 500 -6495 520
rect -4355 500 -4335 520
rect -1475 500 -1455 520
rect -11375 460 -11355 480
rect -6380 460 -6360 480
rect -6200 460 -6180 480
rect -6020 460 -6000 480
rect -5840 460 -5820 480
rect -5660 460 -5640 480
rect -5480 460 -5460 480
rect -5300 460 -5280 480
rect -5120 460 -5100 480
rect -4940 460 -4920 480
rect -4760 460 -4740 480
rect -4580 460 -4560 480
rect -4400 460 -4380 480
rect -11285 420 -11265 440
rect -9980 420 -9960 440
rect -9800 420 -9780 440
rect -9620 420 -9600 440
rect -9440 420 -9420 440
rect -9260 420 -9240 440
rect -9080 420 -9060 440
rect -8900 420 -8880 440
rect -8720 420 -8700 440
rect -8540 420 -8520 440
rect -8360 420 -8340 440
rect -8180 420 -8160 440
rect -8000 420 -7980 440
rect -11195 380 -11175 400
rect -6875 380 -6855 400
rect -6425 380 -6405 400
rect -6245 380 -6225 400
rect -6065 380 -6045 400
rect -5885 380 -5865 400
rect -5705 380 -5685 400
rect -5525 380 -5505 400
rect -5345 380 -5325 400
rect -5165 380 -5145 400
rect -4985 380 -4965 400
rect -4805 380 -4785 400
rect -4625 380 -4605 400
rect -4445 380 -4425 400
rect -3995 380 -3975 400
rect -1835 380 -1815 400
rect -1115 380 -1095 400
rect -11105 340 -11085 360
rect -10475 340 -10455 360
rect -10025 340 -10005 360
rect -9845 340 -9825 360
rect -9665 340 -9645 360
rect -9485 340 -9465 360
rect -9305 340 -9285 360
rect -9125 340 -9105 360
rect -8945 340 -8925 360
rect -8765 340 -8745 360
rect -8585 340 -8565 360
rect -8405 340 -8385 360
rect -8225 340 -8205 360
rect -8045 340 -8025 360
rect -7595 340 -7575 360
rect -3275 340 -3255 360
rect -2555 340 -2535 360
rect -10430 300 -10410 320
rect -10250 300 -10230 320
rect -7910 300 -7890 320
rect -7730 300 -7710 320
rect -6830 300 -6810 320
rect -6650 300 -6630 320
rect -4310 300 -4290 320
rect -4130 300 -4110 320
rect -3230 300 -3210 320
rect -3050 300 -3030 320
rect -2870 300 -2850 320
rect -2690 300 -2670 320
rect -1790 300 -1770 320
rect -1610 300 -1590 320
rect -1430 300 -1410 320
rect -1250 300 -1230 320
rect -215 300 -195 320
rect -10790 260 -10770 280
rect -10610 260 -10590 280
rect -7550 260 -7530 280
rect -7370 260 -7350 280
rect -7190 260 -7170 280
rect -7010 260 -6990 280
rect -3950 260 -3930 280
rect -3770 260 -3750 280
rect -3590 260 -3570 280
rect -3410 260 -3390 280
rect -2510 260 -2490 280
rect -2330 260 -2310 280
rect -2150 260 -2130 280
rect -1970 260 -1950 280
rect -1070 260 -1050 280
rect -890 260 -870 280
rect -125 260 -105 280
rect -10790 175 -10770 195
rect -10610 175 -10590 195
rect -10430 175 -10410 195
rect -10250 175 -10230 195
rect -10070 175 -10050 195
rect -9890 175 -9870 195
rect -9710 175 -9690 195
rect -9530 175 -9510 195
rect -9350 175 -9330 195
rect -9170 175 -9150 195
rect -8990 175 -8970 195
rect -8810 175 -8790 195
rect -8630 175 -8610 195
rect -8450 175 -8430 195
rect -8270 175 -8250 195
rect -8090 175 -8070 195
rect -7910 175 -7890 195
rect -7730 175 -7710 195
rect -7550 175 -7530 195
rect -7370 175 -7350 195
rect -7190 175 -7170 195
rect -7010 175 -6990 195
rect -6830 175 -6810 195
rect -6650 175 -6630 195
rect -6470 175 -6450 195
rect -6290 175 -6270 195
rect -6110 175 -6090 195
rect -5930 175 -5910 195
rect -5750 175 -5730 195
rect -5570 175 -5550 195
rect -5390 175 -5370 195
rect -5210 175 -5190 195
rect -5030 175 -5010 195
rect -4850 175 -4830 195
rect -4670 175 -4650 195
rect -4490 175 -4470 195
rect -4310 175 -4290 195
rect -4130 175 -4110 195
rect -3950 175 -3930 195
rect -3770 175 -3750 195
rect -3590 175 -3570 195
rect -3410 175 -3390 195
rect -3230 175 -3210 195
rect -3050 175 -3030 195
rect -2870 175 -2850 195
rect -2690 175 -2670 195
rect -2510 175 -2490 195
rect -2330 175 -2310 195
rect -2150 175 -2130 195
rect -1970 175 -1950 195
rect -1790 175 -1770 195
rect -1610 175 -1590 195
rect -1430 175 -1410 195
rect -1250 175 -1230 195
rect -1070 175 -1050 195
rect -890 175 -870 195
rect -11555 60 -11535 140
rect -10835 60 -10815 140
rect -10745 60 -10725 140
rect -10655 60 -10635 140
rect -10565 60 -10545 140
rect -10475 60 -10455 140
rect -10385 60 -10365 140
rect -10295 60 -10275 140
rect -10205 60 -10185 140
rect -10115 60 -10095 140
rect -10025 60 -10005 140
rect -9935 60 -9915 140
rect -9845 60 -9825 140
rect -9755 60 -9735 140
rect -9665 60 -9645 140
rect -9575 60 -9555 140
rect -9485 60 -9465 140
rect -9395 60 -9375 140
rect -9305 60 -9285 140
rect -9215 60 -9195 140
rect -9125 60 -9105 140
rect -9035 60 -9015 140
rect -8945 60 -8925 140
rect -8855 60 -8835 140
rect -8765 60 -8745 140
rect -8675 60 -8655 140
rect -8585 60 -8565 140
rect -8495 60 -8475 140
rect -8405 60 -8385 140
rect -8315 60 -8295 140
rect -8225 60 -8205 140
rect -8135 60 -8115 140
rect -8045 60 -8025 140
rect -7955 60 -7935 140
rect -7865 60 -7845 140
rect -7775 60 -7755 140
rect -7685 60 -7665 140
rect -7595 60 -7575 140
rect -7505 60 -7485 140
rect -7415 60 -7395 140
rect -7325 60 -7305 140
rect -7235 60 -7215 140
rect -7145 60 -7125 140
rect -7055 60 -7035 140
rect -6965 60 -6945 140
rect -6875 60 -6855 140
rect -6785 60 -6765 140
rect -6695 60 -6675 140
rect -6605 60 -6585 140
rect -6515 60 -6495 140
rect -6425 60 -6405 140
rect -6335 60 -6315 140
rect -6245 60 -6225 140
rect -6155 60 -6135 140
rect -6065 60 -6045 140
rect -5975 60 -5955 140
rect -5885 60 -5865 140
rect -5795 60 -5775 140
rect -5705 60 -5685 140
rect -5615 60 -5595 140
rect -5525 60 -5505 140
rect -5435 60 -5415 140
rect -5345 60 -5325 140
rect -5255 60 -5235 140
rect -5165 60 -5145 140
rect -5075 60 -5055 140
rect -4985 60 -4965 140
rect -4895 60 -4875 140
rect -4805 60 -4785 140
rect -4715 60 -4695 140
rect -4625 60 -4605 140
rect -4535 60 -4515 140
rect -4445 60 -4425 140
rect -4355 60 -4335 140
rect -4265 60 -4245 140
rect -4175 60 -4155 140
rect -4085 60 -4065 140
rect -3995 60 -3975 140
rect -3905 60 -3885 140
rect -3815 60 -3795 140
rect -3725 60 -3705 140
rect -3635 60 -3615 140
rect -3545 60 -3525 140
rect -3455 60 -3435 140
rect -3365 60 -3345 140
rect -3275 60 -3255 140
rect -3185 60 -3165 140
rect -3095 60 -3075 140
rect -3005 60 -2985 140
rect -2915 60 -2895 140
rect -2825 60 -2805 140
rect -2735 60 -2715 140
rect -2645 60 -2625 140
rect -2555 60 -2535 140
rect -2465 60 -2445 140
rect -2375 60 -2355 140
rect -2285 60 -2265 140
rect -2195 60 -2175 140
rect -2105 60 -2085 140
rect -2015 60 -1995 140
rect -1925 60 -1905 140
rect -1835 60 -1815 140
rect -1745 60 -1725 140
rect -1655 60 -1635 140
rect -1565 60 -1545 140
rect -1475 60 -1455 140
rect -1385 60 -1365 140
rect -1295 60 -1275 140
rect -1205 60 -1185 140
rect -1115 60 -1095 140
rect -1025 60 -1005 140
rect -935 60 -915 140
rect -845 60 -825 140
rect -755 60 -735 140
rect -35 60 -15 140
rect -11690 0 -11670 20
rect -11555 0 -11535 20
rect -10835 0 -10815 20
rect -10655 0 -10635 20
rect -10475 0 -10455 20
rect -10295 0 -10275 20
rect -10115 0 -10095 20
rect -9935 0 -9915 20
rect -9755 0 -9735 20
rect -9575 0 -9555 20
rect -9395 0 -9375 20
rect -9215 0 -9195 20
rect -9035 0 -9015 20
rect -8855 0 -8835 20
rect -8675 0 -8655 20
rect -8495 0 -8475 20
rect -8315 0 -8295 20
rect -8135 0 -8115 20
rect -7955 0 -7935 20
rect -7775 0 -7755 20
rect -7595 0 -7575 20
rect -7415 0 -7395 20
rect -7235 0 -7215 20
rect -7055 0 -7035 20
rect -6875 0 -6855 20
rect -6695 0 -6675 20
rect -6515 0 -6495 20
rect -6335 0 -6315 20
rect -6155 0 -6135 20
rect -5975 0 -5955 20
rect -5795 0 -5775 20
rect -5615 0 -5595 20
rect -5435 0 -5415 20
rect -5255 0 -5235 20
rect -5075 0 -5055 20
rect -4895 0 -4875 20
rect -4715 0 -4695 20
rect -4535 0 -4515 20
rect -4355 0 -4335 20
rect -4175 0 -4155 20
rect -3995 0 -3975 20
rect -3815 0 -3795 20
rect -3635 0 -3615 20
rect -3455 0 -3435 20
rect -3275 0 -3255 20
rect -3095 0 -3075 20
rect -2915 0 -2895 20
rect -2735 0 -2715 20
rect -2555 0 -2535 20
rect -2375 0 -2355 20
rect -2195 0 -2175 20
rect -2015 0 -1995 20
rect -1835 0 -1815 20
rect -1655 0 -1635 20
rect -1475 0 -1455 20
rect -1295 0 -1275 20
rect -1115 0 -1095 20
rect -935 0 -915 20
rect -755 0 -735 20
rect -35 0 -15 20
rect 100 0 120 20
<< metal1 >>
rect -11700 2000 -11660 2005
rect -11700 1970 -11695 2000
rect -11665 1970 -11660 2000
rect -11700 25 -11660 1970
rect -11565 2000 -11525 2005
rect -11565 1970 -11560 2000
rect -11530 1970 -11525 2000
rect -11565 1965 -11525 1970
rect -10845 2000 -10805 2005
rect -10845 1970 -10840 2000
rect -10810 1970 -10805 2000
rect -10845 1965 -10805 1970
rect -10665 2000 -10625 2005
rect -10665 1970 -10660 2000
rect -10630 1970 -10625 2000
rect -10665 1965 -10625 1970
rect -10485 2000 -10445 2005
rect -10485 1970 -10480 2000
rect -10450 1970 -10445 2000
rect -10485 1965 -10445 1970
rect -10305 2000 -10265 2005
rect -10305 1970 -10300 2000
rect -10270 1970 -10265 2000
rect -10305 1965 -10265 1970
rect -10125 2000 -10085 2005
rect -10125 1970 -10120 2000
rect -10090 1970 -10085 2000
rect -10125 1965 -10085 1970
rect -9945 2000 -9905 2005
rect -9945 1970 -9940 2000
rect -9910 1970 -9905 2000
rect -9945 1965 -9905 1970
rect -9765 2000 -9725 2005
rect -9765 1970 -9760 2000
rect -9730 1970 -9725 2000
rect -9765 1965 -9725 1970
rect -9585 2000 -9545 2005
rect -9585 1970 -9580 2000
rect -9550 1970 -9545 2000
rect -9585 1965 -9545 1970
rect -9405 2000 -9365 2005
rect -9405 1970 -9400 2000
rect -9370 1970 -9365 2000
rect -9405 1965 -9365 1970
rect -9225 2000 -9185 2005
rect -9225 1970 -9220 2000
rect -9190 1970 -9185 2000
rect -9225 1965 -9185 1970
rect -9045 2000 -9005 2005
rect -9045 1970 -9040 2000
rect -9010 1970 -9005 2000
rect -9045 1965 -9005 1970
rect -8865 2000 -8825 2005
rect -8865 1970 -8860 2000
rect -8830 1970 -8825 2000
rect -8865 1965 -8825 1970
rect -8685 2000 -8645 2005
rect -8685 1970 -8680 2000
rect -8650 1970 -8645 2000
rect -8685 1965 -8645 1970
rect -8505 2000 -8465 2005
rect -8505 1970 -8500 2000
rect -8470 1970 -8465 2000
rect -8505 1965 -8465 1970
rect -8325 2000 -8285 2005
rect -8325 1970 -8320 2000
rect -8290 1970 -8285 2000
rect -8325 1965 -8285 1970
rect -8145 2000 -8105 2005
rect -8145 1970 -8140 2000
rect -8110 1970 -8105 2000
rect -8145 1965 -8105 1970
rect -7965 2000 -7925 2005
rect -7965 1970 -7960 2000
rect -7930 1970 -7925 2000
rect -7965 1965 -7925 1970
rect -7785 2000 -7745 2005
rect -7785 1970 -7780 2000
rect -7750 1970 -7745 2000
rect -7785 1965 -7745 1970
rect -7605 2000 -7565 2005
rect -7605 1970 -7600 2000
rect -7570 1970 -7565 2000
rect -7605 1965 -7565 1970
rect -7425 2000 -7385 2005
rect -7425 1970 -7420 2000
rect -7390 1970 -7385 2000
rect -7425 1965 -7385 1970
rect -7245 2000 -7205 2005
rect -7245 1970 -7240 2000
rect -7210 1970 -7205 2000
rect -7245 1965 -7205 1970
rect -7065 2000 -7025 2005
rect -7065 1970 -7060 2000
rect -7030 1970 -7025 2000
rect -7065 1965 -7025 1970
rect -6885 2000 -6845 2005
rect -6885 1970 -6880 2000
rect -6850 1970 -6845 2000
rect -6885 1965 -6845 1970
rect -6705 2000 -6665 2005
rect -6705 1970 -6700 2000
rect -6670 1970 -6665 2000
rect -6705 1965 -6665 1970
rect -6525 2000 -6485 2005
rect -6525 1970 -6520 2000
rect -6490 1970 -6485 2000
rect -6525 1965 -6485 1970
rect -6345 2000 -6305 2005
rect -6345 1970 -6340 2000
rect -6310 1970 -6305 2000
rect -6345 1965 -6305 1970
rect -6165 2000 -6125 2005
rect -6165 1970 -6160 2000
rect -6130 1970 -6125 2000
rect -6165 1965 -6125 1970
rect -5985 2000 -5945 2005
rect -5985 1970 -5980 2000
rect -5950 1970 -5945 2000
rect -5985 1965 -5945 1970
rect -5805 2000 -5765 2005
rect -5805 1970 -5800 2000
rect -5770 1970 -5765 2000
rect -5805 1965 -5765 1970
rect -5625 2000 -5585 2005
rect -5625 1970 -5620 2000
rect -5590 1970 -5585 2000
rect -5625 1965 -5585 1970
rect -5445 2000 -5405 2005
rect -5445 1970 -5440 2000
rect -5410 1970 -5405 2000
rect -5445 1965 -5405 1970
rect -5265 2000 -5225 2005
rect -5265 1970 -5260 2000
rect -5230 1970 -5225 2000
rect -5265 1965 -5225 1970
rect -5085 2000 -5045 2005
rect -5085 1970 -5080 2000
rect -5050 1970 -5045 2000
rect -5085 1965 -5045 1970
rect -4905 2000 -4865 2005
rect -4905 1970 -4900 2000
rect -4870 1970 -4865 2000
rect -4905 1965 -4865 1970
rect -4725 2000 -4685 2005
rect -4725 1970 -4720 2000
rect -4690 1970 -4685 2000
rect -4725 1965 -4685 1970
rect -4545 2000 -4505 2005
rect -4545 1970 -4540 2000
rect -4510 1970 -4505 2000
rect -4545 1965 -4505 1970
rect -4365 2000 -4325 2005
rect -4365 1970 -4360 2000
rect -4330 1970 -4325 2000
rect -4365 1965 -4325 1970
rect -4185 2000 -4145 2005
rect -4185 1970 -4180 2000
rect -4150 1970 -4145 2000
rect -4185 1965 -4145 1970
rect -4005 2000 -3965 2005
rect -4005 1970 -4000 2000
rect -3970 1970 -3965 2000
rect -4005 1965 -3965 1970
rect -3825 2000 -3785 2005
rect -3825 1970 -3820 2000
rect -3790 1970 -3785 2000
rect -3825 1965 -3785 1970
rect -3645 2000 -3605 2005
rect -3645 1970 -3640 2000
rect -3610 1970 -3605 2000
rect -3645 1965 -3605 1970
rect -3465 2000 -3425 2005
rect -3465 1970 -3460 2000
rect -3430 1970 -3425 2000
rect -3465 1965 -3425 1970
rect -3285 2000 -3245 2005
rect -3285 1970 -3280 2000
rect -3250 1970 -3245 2000
rect -3285 1965 -3245 1970
rect -3105 2000 -3065 2005
rect -3105 1970 -3100 2000
rect -3070 1970 -3065 2000
rect -3105 1965 -3065 1970
rect -2925 2000 -2885 2005
rect -2925 1970 -2920 2000
rect -2890 1970 -2885 2000
rect -2925 1965 -2885 1970
rect -2745 2000 -2705 2005
rect -2745 1970 -2740 2000
rect -2710 1970 -2705 2000
rect -2745 1965 -2705 1970
rect -2565 2000 -2525 2005
rect -2565 1970 -2560 2000
rect -2530 1970 -2525 2000
rect -2565 1965 -2525 1970
rect -2385 2000 -2345 2005
rect -2385 1970 -2380 2000
rect -2350 1970 -2345 2000
rect -2385 1965 -2345 1970
rect -2205 2000 -2165 2005
rect -2205 1970 -2200 2000
rect -2170 1970 -2165 2000
rect -2205 1965 -2165 1970
rect -2025 2000 -1985 2005
rect -2025 1970 -2020 2000
rect -1990 1970 -1985 2000
rect -2025 1965 -1985 1970
rect -1845 2000 -1805 2005
rect -1845 1970 -1840 2000
rect -1810 1970 -1805 2000
rect -1845 1965 -1805 1970
rect -1665 2000 -1625 2005
rect -1665 1970 -1660 2000
rect -1630 1970 -1625 2000
rect -1665 1965 -1625 1970
rect -1485 2000 -1445 2005
rect -1485 1970 -1480 2000
rect -1450 1970 -1445 2000
rect -1485 1965 -1445 1970
rect -1305 2000 -1265 2005
rect -1305 1970 -1300 2000
rect -1270 1970 -1265 2000
rect -1305 1965 -1265 1970
rect -1125 2000 -1085 2005
rect -1125 1970 -1120 2000
rect -1090 1970 -1085 2000
rect -1125 1965 -1085 1970
rect -945 2000 -905 2005
rect -945 1970 -940 2000
rect -910 1970 -905 2000
rect -945 1965 -905 1970
rect -765 2000 -725 2005
rect -765 1970 -760 2000
rect -730 1970 -725 2000
rect -765 1965 -725 1970
rect -45 2000 -5 2005
rect -45 1970 -40 2000
rect -10 1970 -5 2000
rect -45 1965 -5 1970
rect 90 2000 130 2005
rect 90 1970 95 2000
rect 125 1970 130 2000
rect -11555 1945 -11535 1965
rect -10835 1945 -10815 1965
rect -9395 1945 -9375 1965
rect -7955 1945 -7935 1965
rect -4355 1945 -4335 1965
rect -755 1945 -735 1965
rect -35 1945 -15 1965
rect -11560 1935 -11530 1945
rect -11560 1855 -11555 1935
rect -11535 1855 -11530 1935
rect -11560 1845 -11530 1855
rect -11470 1845 -11440 1945
rect -11380 1845 -11350 1945
rect -11290 1845 -11260 1945
rect -11200 1845 -11170 1945
rect -11110 1845 -11080 1945
rect -11020 1845 -10990 1945
rect -10930 1845 -10900 1945
rect -10840 1935 -10810 1945
rect -10840 1855 -10835 1935
rect -10815 1855 -10810 1935
rect -10840 1845 -10810 1855
rect -10750 1935 -10720 1945
rect -10750 1855 -10745 1935
rect -10725 1855 -10720 1935
rect -10750 1845 -10720 1855
rect -10660 1935 -10630 1945
rect -10660 1855 -10655 1935
rect -10635 1855 -10630 1935
rect -10660 1845 -10630 1855
rect -10570 1935 -10540 1945
rect -10570 1855 -10565 1935
rect -10545 1855 -10540 1935
rect -10570 1845 -10540 1855
rect -10480 1935 -10450 1945
rect -10480 1855 -10475 1935
rect -10455 1855 -10450 1935
rect -10480 1845 -10450 1855
rect -10390 1935 -10360 1945
rect -10390 1855 -10385 1935
rect -10365 1855 -10360 1935
rect -10390 1845 -10360 1855
rect -10300 1935 -10270 1945
rect -10300 1855 -10295 1935
rect -10275 1855 -10270 1935
rect -10300 1845 -10270 1855
rect -10210 1935 -10180 1945
rect -10210 1855 -10205 1935
rect -10185 1855 -10180 1935
rect -10210 1845 -10180 1855
rect -10120 1935 -10090 1945
rect -10120 1855 -10115 1935
rect -10095 1855 -10090 1935
rect -10120 1845 -10090 1855
rect -10030 1935 -10000 1945
rect -10030 1855 -10025 1935
rect -10005 1855 -10000 1935
rect -10030 1845 -10000 1855
rect -9940 1935 -9910 1945
rect -9940 1855 -9935 1935
rect -9915 1855 -9910 1935
rect -9940 1845 -9910 1855
rect -9850 1935 -9820 1945
rect -9850 1855 -9845 1935
rect -9825 1855 -9820 1935
rect -9850 1845 -9820 1855
rect -9760 1935 -9730 1945
rect -9760 1855 -9755 1935
rect -9735 1855 -9730 1935
rect -9760 1845 -9730 1855
rect -9670 1935 -9640 1945
rect -9670 1855 -9665 1935
rect -9645 1855 -9640 1935
rect -9670 1845 -9640 1855
rect -9580 1935 -9550 1945
rect -9580 1855 -9575 1935
rect -9555 1855 -9550 1935
rect -9580 1845 -9550 1855
rect -9490 1935 -9460 1945
rect -9490 1855 -9485 1935
rect -9465 1855 -9460 1935
rect -9490 1845 -9460 1855
rect -9400 1935 -9370 1945
rect -9400 1855 -9395 1935
rect -9375 1855 -9370 1935
rect -9400 1845 -9370 1855
rect -9310 1935 -9280 1945
rect -9310 1855 -9305 1935
rect -9285 1855 -9280 1935
rect -9310 1845 -9280 1855
rect -9220 1935 -9190 1945
rect -9220 1855 -9215 1935
rect -9195 1855 -9190 1935
rect -9220 1845 -9190 1855
rect -9130 1935 -9100 1945
rect -9130 1855 -9125 1935
rect -9105 1855 -9100 1935
rect -9130 1845 -9100 1855
rect -9040 1935 -9010 1945
rect -9040 1855 -9035 1935
rect -9015 1855 -9010 1935
rect -9040 1845 -9010 1855
rect -8950 1935 -8920 1945
rect -8950 1855 -8945 1935
rect -8925 1855 -8920 1935
rect -8950 1845 -8920 1855
rect -8860 1935 -8830 1945
rect -8860 1855 -8855 1935
rect -8835 1855 -8830 1935
rect -8860 1845 -8830 1855
rect -8770 1935 -8740 1945
rect -8770 1855 -8765 1935
rect -8745 1855 -8740 1935
rect -8770 1845 -8740 1855
rect -8680 1935 -8650 1945
rect -8680 1855 -8675 1935
rect -8655 1855 -8650 1935
rect -8680 1845 -8650 1855
rect -8590 1935 -8560 1945
rect -8590 1855 -8585 1935
rect -8565 1855 -8560 1935
rect -8590 1845 -8560 1855
rect -8500 1935 -8470 1945
rect -8500 1855 -8495 1935
rect -8475 1855 -8470 1935
rect -8500 1845 -8470 1855
rect -8410 1935 -8380 1945
rect -8410 1855 -8405 1935
rect -8385 1855 -8380 1935
rect -8410 1845 -8380 1855
rect -8320 1935 -8290 1945
rect -8320 1855 -8315 1935
rect -8295 1855 -8290 1935
rect -8320 1845 -8290 1855
rect -8230 1935 -8200 1945
rect -8230 1855 -8225 1935
rect -8205 1855 -8200 1935
rect -8230 1845 -8200 1855
rect -8140 1935 -8110 1945
rect -8140 1855 -8135 1935
rect -8115 1855 -8110 1935
rect -8140 1845 -8110 1855
rect -8050 1935 -8020 1945
rect -8050 1855 -8045 1935
rect -8025 1855 -8020 1935
rect -8050 1845 -8020 1855
rect -7960 1935 -7930 1945
rect -7960 1855 -7955 1935
rect -7935 1855 -7930 1935
rect -7960 1845 -7930 1855
rect -7870 1935 -7840 1945
rect -7870 1855 -7865 1935
rect -7845 1855 -7840 1935
rect -7870 1845 -7840 1855
rect -7780 1935 -7750 1945
rect -7780 1855 -7775 1935
rect -7755 1855 -7750 1935
rect -7780 1845 -7750 1855
rect -7690 1935 -7660 1945
rect -7690 1855 -7685 1935
rect -7665 1855 -7660 1935
rect -7690 1845 -7660 1855
rect -7600 1935 -7570 1945
rect -7600 1855 -7595 1935
rect -7575 1855 -7570 1935
rect -7600 1845 -7570 1855
rect -7510 1935 -7480 1945
rect -7510 1855 -7505 1935
rect -7485 1855 -7480 1935
rect -7510 1845 -7480 1855
rect -7420 1935 -7390 1945
rect -7420 1855 -7415 1935
rect -7395 1855 -7390 1935
rect -7420 1845 -7390 1855
rect -7330 1935 -7300 1945
rect -7330 1855 -7325 1935
rect -7305 1855 -7300 1935
rect -7330 1845 -7300 1855
rect -7240 1935 -7210 1945
rect -7240 1855 -7235 1935
rect -7215 1855 -7210 1935
rect -7240 1845 -7210 1855
rect -7150 1935 -7120 1945
rect -7150 1855 -7145 1935
rect -7125 1855 -7120 1935
rect -7150 1845 -7120 1855
rect -7060 1935 -7030 1945
rect -7060 1855 -7055 1935
rect -7035 1855 -7030 1935
rect -7060 1845 -7030 1855
rect -6970 1935 -6940 1945
rect -6970 1855 -6965 1935
rect -6945 1855 -6940 1935
rect -6970 1845 -6940 1855
rect -6880 1935 -6850 1945
rect -6880 1855 -6875 1935
rect -6855 1855 -6850 1935
rect -6880 1845 -6850 1855
rect -6790 1935 -6760 1945
rect -6790 1855 -6785 1935
rect -6765 1855 -6760 1935
rect -6790 1845 -6760 1855
rect -6700 1935 -6670 1945
rect -6700 1855 -6695 1935
rect -6675 1855 -6670 1935
rect -6700 1845 -6670 1855
rect -6610 1935 -6580 1945
rect -6610 1855 -6605 1935
rect -6585 1855 -6580 1935
rect -6610 1845 -6580 1855
rect -6520 1935 -6490 1945
rect -6520 1855 -6515 1935
rect -6495 1855 -6490 1935
rect -6520 1845 -6490 1855
rect -6430 1935 -6400 1945
rect -6430 1855 -6425 1935
rect -6405 1855 -6400 1935
rect -6430 1845 -6400 1855
rect -6340 1935 -6310 1945
rect -6340 1855 -6335 1935
rect -6315 1855 -6310 1935
rect -6340 1845 -6310 1855
rect -6250 1935 -6220 1945
rect -6250 1855 -6245 1935
rect -6225 1855 -6220 1935
rect -6250 1845 -6220 1855
rect -6160 1935 -6130 1945
rect -6160 1855 -6155 1935
rect -6135 1855 -6130 1935
rect -6160 1845 -6130 1855
rect -6070 1935 -6040 1945
rect -6070 1855 -6065 1935
rect -6045 1855 -6040 1935
rect -6070 1845 -6040 1855
rect -5980 1935 -5950 1945
rect -5980 1855 -5975 1935
rect -5955 1855 -5950 1935
rect -5980 1845 -5950 1855
rect -5890 1935 -5860 1945
rect -5890 1855 -5885 1935
rect -5865 1855 -5860 1935
rect -5890 1845 -5860 1855
rect -5800 1935 -5770 1945
rect -5800 1855 -5795 1935
rect -5775 1855 -5770 1935
rect -5800 1845 -5770 1855
rect -5710 1935 -5680 1945
rect -5710 1855 -5705 1935
rect -5685 1855 -5680 1935
rect -5710 1845 -5680 1855
rect -5620 1935 -5590 1945
rect -5620 1855 -5615 1935
rect -5595 1855 -5590 1935
rect -5620 1845 -5590 1855
rect -5530 1935 -5500 1945
rect -5530 1855 -5525 1935
rect -5505 1855 -5500 1935
rect -5530 1845 -5500 1855
rect -5440 1935 -5410 1945
rect -5440 1855 -5435 1935
rect -5415 1855 -5410 1935
rect -5440 1845 -5410 1855
rect -5350 1935 -5320 1945
rect -5350 1855 -5345 1935
rect -5325 1855 -5320 1935
rect -5350 1845 -5320 1855
rect -5260 1935 -5230 1945
rect -5260 1855 -5255 1935
rect -5235 1855 -5230 1935
rect -5260 1845 -5230 1855
rect -5170 1935 -5140 1945
rect -5170 1855 -5165 1935
rect -5145 1855 -5140 1935
rect -5170 1845 -5140 1855
rect -5080 1935 -5050 1945
rect -5080 1855 -5075 1935
rect -5055 1855 -5050 1935
rect -5080 1845 -5050 1855
rect -4990 1935 -4960 1945
rect -4990 1855 -4985 1935
rect -4965 1855 -4960 1935
rect -4990 1845 -4960 1855
rect -4900 1935 -4870 1945
rect -4900 1855 -4895 1935
rect -4875 1855 -4870 1935
rect -4900 1845 -4870 1855
rect -4810 1935 -4780 1945
rect -4810 1855 -4805 1935
rect -4785 1855 -4780 1935
rect -4810 1845 -4780 1855
rect -4720 1935 -4690 1945
rect -4720 1855 -4715 1935
rect -4695 1855 -4690 1935
rect -4720 1845 -4690 1855
rect -4630 1935 -4600 1945
rect -4630 1855 -4625 1935
rect -4605 1855 -4600 1935
rect -4630 1845 -4600 1855
rect -4540 1935 -4510 1945
rect -4540 1855 -4535 1935
rect -4515 1855 -4510 1935
rect -4540 1845 -4510 1855
rect -4450 1935 -4420 1945
rect -4450 1855 -4445 1935
rect -4425 1855 -4420 1935
rect -4450 1845 -4420 1855
rect -4360 1935 -4330 1945
rect -4360 1855 -4355 1935
rect -4335 1855 -4330 1935
rect -4360 1845 -4330 1855
rect -4270 1935 -4240 1945
rect -4270 1855 -4265 1935
rect -4245 1855 -4240 1935
rect -4270 1845 -4240 1855
rect -4180 1935 -4150 1945
rect -4180 1855 -4175 1935
rect -4155 1855 -4150 1935
rect -4180 1845 -4150 1855
rect -4090 1935 -4060 1945
rect -4090 1855 -4085 1935
rect -4065 1855 -4060 1935
rect -4090 1845 -4060 1855
rect -4000 1935 -3970 1945
rect -4000 1855 -3995 1935
rect -3975 1855 -3970 1935
rect -4000 1845 -3970 1855
rect -3910 1935 -3880 1945
rect -3910 1855 -3905 1935
rect -3885 1855 -3880 1935
rect -3910 1845 -3880 1855
rect -3820 1935 -3790 1945
rect -3820 1855 -3815 1935
rect -3795 1855 -3790 1935
rect -3820 1845 -3790 1855
rect -3730 1935 -3700 1945
rect -3730 1855 -3725 1935
rect -3705 1855 -3700 1935
rect -3730 1845 -3700 1855
rect -3640 1935 -3610 1945
rect -3640 1855 -3635 1935
rect -3615 1855 -3610 1935
rect -3640 1845 -3610 1855
rect -3550 1935 -3520 1945
rect -3550 1855 -3545 1935
rect -3525 1855 -3520 1935
rect -3550 1845 -3520 1855
rect -3460 1935 -3430 1945
rect -3460 1855 -3455 1935
rect -3435 1855 -3430 1935
rect -3460 1845 -3430 1855
rect -3370 1935 -3340 1945
rect -3370 1855 -3365 1935
rect -3345 1855 -3340 1935
rect -3370 1845 -3340 1855
rect -3280 1935 -3250 1945
rect -3280 1855 -3275 1935
rect -3255 1855 -3250 1935
rect -3280 1845 -3250 1855
rect -3190 1935 -3160 1945
rect -3190 1855 -3185 1935
rect -3165 1855 -3160 1935
rect -3190 1845 -3160 1855
rect -3100 1935 -3070 1945
rect -3100 1855 -3095 1935
rect -3075 1855 -3070 1935
rect -3100 1845 -3070 1855
rect -3010 1935 -2980 1945
rect -3010 1855 -3005 1935
rect -2985 1855 -2980 1935
rect -3010 1845 -2980 1855
rect -2920 1935 -2890 1945
rect -2920 1855 -2915 1935
rect -2895 1855 -2890 1935
rect -2920 1845 -2890 1855
rect -2830 1935 -2800 1945
rect -2830 1855 -2825 1935
rect -2805 1855 -2800 1935
rect -2830 1845 -2800 1855
rect -2740 1935 -2710 1945
rect -2740 1855 -2735 1935
rect -2715 1855 -2710 1935
rect -2740 1845 -2710 1855
rect -2650 1935 -2620 1945
rect -2650 1855 -2645 1935
rect -2625 1855 -2620 1935
rect -2650 1845 -2620 1855
rect -2560 1935 -2530 1945
rect -2560 1855 -2555 1935
rect -2535 1855 -2530 1935
rect -2560 1845 -2530 1855
rect -2470 1935 -2440 1945
rect -2470 1855 -2465 1935
rect -2445 1855 -2440 1935
rect -2470 1845 -2440 1855
rect -2380 1935 -2350 1945
rect -2380 1855 -2375 1935
rect -2355 1855 -2350 1935
rect -2380 1845 -2350 1855
rect -2290 1935 -2260 1945
rect -2290 1855 -2285 1935
rect -2265 1855 -2260 1935
rect -2290 1845 -2260 1855
rect -2200 1935 -2170 1945
rect -2200 1855 -2195 1935
rect -2175 1855 -2170 1935
rect -2200 1845 -2170 1855
rect -2110 1935 -2080 1945
rect -2110 1855 -2105 1935
rect -2085 1855 -2080 1935
rect -2110 1845 -2080 1855
rect -2020 1935 -1990 1945
rect -2020 1855 -2015 1935
rect -1995 1855 -1990 1935
rect -2020 1845 -1990 1855
rect -1930 1935 -1900 1945
rect -1930 1855 -1925 1935
rect -1905 1855 -1900 1935
rect -1930 1845 -1900 1855
rect -1840 1935 -1810 1945
rect -1840 1855 -1835 1935
rect -1815 1855 -1810 1935
rect -1840 1845 -1810 1855
rect -1750 1935 -1720 1945
rect -1750 1855 -1745 1935
rect -1725 1855 -1720 1935
rect -1750 1845 -1720 1855
rect -1660 1935 -1630 1945
rect -1660 1855 -1655 1935
rect -1635 1855 -1630 1935
rect -1660 1845 -1630 1855
rect -1570 1935 -1540 1945
rect -1570 1855 -1565 1935
rect -1545 1855 -1540 1935
rect -1570 1845 -1540 1855
rect -1480 1935 -1450 1945
rect -1480 1855 -1475 1935
rect -1455 1855 -1450 1935
rect -1480 1845 -1450 1855
rect -1390 1935 -1360 1945
rect -1390 1855 -1385 1935
rect -1365 1855 -1360 1935
rect -1390 1845 -1360 1855
rect -1300 1935 -1270 1945
rect -1300 1855 -1295 1935
rect -1275 1855 -1270 1935
rect -1300 1845 -1270 1855
rect -1210 1935 -1180 1945
rect -1210 1855 -1205 1935
rect -1185 1855 -1180 1935
rect -1210 1845 -1180 1855
rect -1120 1935 -1090 1945
rect -1120 1855 -1115 1935
rect -1095 1855 -1090 1935
rect -1120 1845 -1090 1855
rect -1030 1935 -1000 1945
rect -1030 1855 -1025 1935
rect -1005 1855 -1000 1935
rect -1030 1845 -1000 1855
rect -940 1935 -910 1945
rect -940 1855 -935 1935
rect -915 1855 -910 1935
rect -940 1845 -910 1855
rect -850 1935 -820 1945
rect -850 1855 -845 1935
rect -825 1855 -820 1935
rect -850 1845 -820 1855
rect -760 1935 -730 1945
rect -760 1855 -755 1935
rect -735 1855 -730 1935
rect -760 1845 -730 1855
rect -670 1845 -640 1945
rect -580 1845 -550 1945
rect -490 1845 -460 1945
rect -400 1845 -370 1945
rect -310 1845 -280 1945
rect -220 1845 -190 1945
rect -130 1845 -100 1945
rect -40 1935 -10 1945
rect -40 1855 -35 1935
rect -15 1855 -10 1935
rect -40 1845 -10 1855
rect -11465 1500 -11445 1845
rect -11375 1540 -11355 1845
rect -11285 1580 -11265 1845
rect -11195 1620 -11175 1845
rect -11105 1660 -11085 1845
rect -11110 1655 -11080 1660
rect -11110 1635 -11105 1655
rect -11085 1635 -11080 1655
rect -11110 1630 -11080 1635
rect -11200 1615 -11170 1620
rect -11200 1595 -11195 1615
rect -11175 1595 -11170 1615
rect -11200 1590 -11170 1595
rect -11290 1575 -11260 1580
rect -11290 1555 -11285 1575
rect -11265 1555 -11260 1575
rect -11290 1550 -11260 1555
rect -11380 1535 -11350 1540
rect -11380 1515 -11375 1535
rect -11355 1515 -11350 1535
rect -11380 1510 -11350 1515
rect -11470 1495 -11440 1500
rect -11470 1475 -11465 1495
rect -11445 1475 -11440 1495
rect -11470 1470 -11440 1475
rect -11465 1165 -11445 1470
rect -11375 1165 -11355 1510
rect -11285 1165 -11265 1550
rect -11195 1165 -11175 1590
rect -11105 1165 -11085 1630
rect -11015 1165 -10995 1845
rect -10925 1165 -10905 1845
rect -10700 1825 -10680 1830
rect -10520 1825 -10500 1830
rect -10705 1820 -10675 1825
rect -10705 1800 -10700 1820
rect -10680 1800 -10675 1820
rect -10705 1795 -10675 1800
rect -10525 1820 -10495 1825
rect -10525 1800 -10520 1820
rect -10500 1800 -10495 1820
rect -10525 1795 -10495 1800
rect -10700 1740 -10680 1795
rect -10520 1740 -10500 1795
rect -10705 1735 -10675 1740
rect -10705 1715 -10700 1735
rect -10680 1715 -10675 1735
rect -10705 1710 -10675 1715
rect -10525 1735 -10495 1740
rect -10525 1715 -10520 1735
rect -10500 1715 -10495 1735
rect -10525 1710 -10495 1715
rect -10700 1705 -10680 1710
rect -10520 1705 -10500 1710
rect -10475 1620 -10455 1845
rect -10340 1825 -10320 1830
rect -10160 1825 -10140 1830
rect -10345 1820 -10315 1825
rect -10345 1800 -10340 1820
rect -10320 1800 -10315 1820
rect -10345 1795 -10315 1800
rect -10165 1820 -10135 1825
rect -10165 1800 -10160 1820
rect -10140 1800 -10135 1820
rect -10165 1795 -10135 1800
rect -10340 1700 -10320 1795
rect -10160 1700 -10140 1795
rect -10345 1695 -10315 1700
rect -10345 1675 -10340 1695
rect -10320 1675 -10315 1695
rect -10345 1670 -10315 1675
rect -10165 1695 -10135 1700
rect -10165 1675 -10160 1695
rect -10140 1675 -10135 1695
rect -10165 1670 -10135 1675
rect -10340 1665 -10320 1670
rect -10160 1665 -10140 1670
rect -10480 1615 -10450 1620
rect -10480 1595 -10475 1615
rect -10455 1595 -10450 1615
rect -10480 1590 -10450 1595
rect -10475 1585 -10455 1590
rect -10115 1500 -10095 1845
rect -9980 1825 -9960 1830
rect -9800 1825 -9780 1830
rect -9985 1820 -9955 1825
rect -9985 1800 -9980 1820
rect -9960 1800 -9955 1820
rect -9985 1795 -9955 1800
rect -9805 1820 -9775 1825
rect -9805 1800 -9800 1820
rect -9780 1800 -9775 1820
rect -9805 1795 -9775 1800
rect -9980 1700 -9960 1795
rect -9800 1700 -9780 1795
rect -9985 1695 -9955 1700
rect -9985 1675 -9980 1695
rect -9960 1675 -9955 1695
rect -9985 1670 -9955 1675
rect -9805 1695 -9775 1700
rect -9805 1675 -9800 1695
rect -9780 1675 -9775 1695
rect -9805 1670 -9775 1675
rect -9980 1665 -9960 1670
rect -9800 1665 -9780 1670
rect -9755 1620 -9735 1845
rect -9620 1825 -9600 1830
rect -9440 1825 -9420 1830
rect -9260 1825 -9240 1830
rect -9080 1825 -9060 1830
rect -9625 1820 -9595 1825
rect -9625 1800 -9620 1820
rect -9600 1800 -9595 1820
rect -9625 1795 -9595 1800
rect -9445 1820 -9415 1825
rect -9445 1800 -9440 1820
rect -9420 1800 -9415 1820
rect -9445 1795 -9415 1800
rect -9265 1820 -9235 1825
rect -9265 1800 -9260 1820
rect -9240 1800 -9235 1820
rect -9265 1795 -9235 1800
rect -9085 1820 -9055 1825
rect -9085 1800 -9080 1820
rect -9060 1800 -9055 1820
rect -9085 1795 -9055 1800
rect -9620 1740 -9600 1795
rect -9440 1740 -9420 1795
rect -9260 1740 -9240 1795
rect -9080 1740 -9060 1795
rect -9625 1735 -9595 1740
rect -9625 1715 -9620 1735
rect -9600 1715 -9595 1735
rect -9625 1710 -9595 1715
rect -9445 1735 -9415 1740
rect -9445 1715 -9440 1735
rect -9420 1715 -9415 1735
rect -9445 1710 -9415 1715
rect -9265 1735 -9235 1740
rect -9265 1715 -9260 1735
rect -9240 1715 -9235 1735
rect -9265 1710 -9235 1715
rect -9085 1735 -9055 1740
rect -9085 1715 -9080 1735
rect -9060 1715 -9055 1735
rect -9085 1710 -9055 1715
rect -9620 1705 -9600 1710
rect -9440 1705 -9420 1710
rect -9260 1705 -9240 1710
rect -9080 1705 -9060 1710
rect -9035 1660 -9015 1845
rect -8900 1825 -8880 1830
rect -8720 1825 -8700 1830
rect -8905 1820 -8875 1825
rect -8905 1800 -8900 1820
rect -8880 1800 -8875 1820
rect -8905 1795 -8875 1800
rect -8725 1820 -8695 1825
rect -8725 1800 -8720 1820
rect -8700 1800 -8695 1820
rect -8725 1795 -8695 1800
rect -8900 1700 -8880 1795
rect -8720 1700 -8700 1795
rect -8905 1695 -8875 1700
rect -8905 1675 -8900 1695
rect -8880 1675 -8875 1695
rect -8905 1670 -8875 1675
rect -8725 1695 -8695 1700
rect -8725 1675 -8720 1695
rect -8700 1675 -8695 1695
rect -8725 1670 -8695 1675
rect -8900 1665 -8880 1670
rect -8720 1665 -8700 1670
rect -9040 1655 -9010 1660
rect -9040 1635 -9035 1655
rect -9015 1635 -9010 1655
rect -9040 1630 -9010 1635
rect -9035 1625 -9015 1630
rect -9760 1615 -9730 1620
rect -9760 1595 -9755 1615
rect -9735 1595 -9730 1615
rect -9760 1590 -9730 1595
rect -9755 1585 -9735 1590
rect -10120 1495 -10090 1500
rect -10120 1475 -10115 1495
rect -10095 1475 -10090 1495
rect -10120 1470 -10090 1475
rect -10790 1460 -10770 1465
rect -10610 1460 -10590 1465
rect -10795 1455 -10765 1460
rect -10795 1435 -10790 1455
rect -10770 1435 -10765 1455
rect -10795 1430 -10765 1435
rect -10615 1455 -10585 1460
rect -10615 1435 -10610 1455
rect -10590 1435 -10585 1455
rect -10615 1430 -10585 1435
rect -10790 1215 -10770 1430
rect -10610 1215 -10590 1430
rect -10430 1420 -10410 1425
rect -10250 1420 -10230 1425
rect -10435 1415 -10405 1420
rect -10435 1395 -10430 1415
rect -10410 1395 -10405 1415
rect -10435 1390 -10405 1395
rect -10255 1415 -10225 1420
rect -10255 1395 -10250 1415
rect -10230 1395 -10225 1415
rect -10255 1390 -10225 1395
rect -10430 1215 -10410 1390
rect -10250 1215 -10230 1390
rect -10795 1210 -10765 1215
rect -10795 1190 -10790 1210
rect -10770 1190 -10765 1210
rect -10795 1185 -10765 1190
rect -10615 1210 -10585 1215
rect -10615 1190 -10610 1210
rect -10590 1190 -10585 1210
rect -10615 1185 -10585 1190
rect -10435 1210 -10405 1215
rect -10435 1190 -10430 1210
rect -10410 1190 -10405 1210
rect -10435 1185 -10405 1190
rect -10255 1210 -10225 1215
rect -10255 1190 -10250 1210
rect -10230 1190 -10225 1210
rect -10255 1185 -10225 1190
rect -10790 1180 -10770 1185
rect -10610 1180 -10590 1185
rect -10430 1180 -10410 1185
rect -10250 1180 -10230 1185
rect -10115 1165 -10095 1470
rect -9710 1460 -9690 1465
rect -9530 1460 -9510 1465
rect -9350 1460 -9330 1465
rect -9170 1460 -9150 1465
rect -8675 1460 -8655 1845
rect -8540 1825 -8520 1830
rect -8360 1825 -8340 1830
rect -8545 1820 -8515 1825
rect -8545 1800 -8540 1820
rect -8520 1800 -8515 1820
rect -8545 1795 -8515 1800
rect -8365 1820 -8335 1825
rect -8365 1800 -8360 1820
rect -8340 1800 -8335 1820
rect -8365 1795 -8335 1800
rect -8540 1700 -8520 1795
rect -8360 1700 -8340 1795
rect -8545 1695 -8515 1700
rect -8545 1675 -8540 1695
rect -8520 1675 -8515 1695
rect -8545 1670 -8515 1675
rect -8365 1695 -8335 1700
rect -8365 1675 -8360 1695
rect -8340 1675 -8335 1695
rect -8365 1670 -8335 1675
rect -8540 1665 -8520 1670
rect -8360 1665 -8340 1670
rect -8315 1660 -8295 1845
rect -8180 1825 -8160 1830
rect -8000 1825 -7980 1830
rect -7820 1825 -7800 1830
rect -7640 1825 -7620 1830
rect -8185 1820 -8155 1825
rect -8185 1800 -8180 1820
rect -8160 1800 -8155 1820
rect -8185 1795 -8155 1800
rect -8005 1820 -7975 1825
rect -8005 1800 -8000 1820
rect -7980 1800 -7975 1820
rect -8005 1795 -7975 1800
rect -7825 1820 -7795 1825
rect -7825 1800 -7820 1820
rect -7800 1800 -7795 1820
rect -7825 1795 -7795 1800
rect -7645 1820 -7615 1825
rect -7645 1800 -7640 1820
rect -7620 1800 -7615 1820
rect -7645 1795 -7615 1800
rect -8180 1740 -8160 1795
rect -8000 1740 -7980 1795
rect -7820 1740 -7800 1795
rect -7640 1740 -7620 1795
rect -8185 1735 -8155 1740
rect -8185 1715 -8180 1735
rect -8160 1715 -8155 1735
rect -8185 1710 -8155 1715
rect -8005 1735 -7975 1740
rect -8005 1715 -8000 1735
rect -7980 1715 -7975 1735
rect -8005 1710 -7975 1715
rect -7825 1735 -7795 1740
rect -7825 1715 -7820 1735
rect -7800 1715 -7795 1735
rect -7825 1710 -7795 1715
rect -7645 1735 -7615 1740
rect -7645 1715 -7640 1735
rect -7620 1715 -7615 1735
rect -7645 1710 -7615 1715
rect -8180 1705 -8160 1710
rect -8000 1705 -7980 1710
rect -7820 1705 -7800 1710
rect -7640 1705 -7620 1710
rect -8320 1655 -8290 1660
rect -8320 1635 -8315 1655
rect -8295 1635 -8290 1655
rect -8320 1630 -8290 1635
rect -8315 1625 -8295 1630
rect -7595 1620 -7575 1845
rect -7460 1825 -7440 1830
rect -7280 1825 -7260 1830
rect -7465 1820 -7435 1825
rect -7465 1800 -7460 1820
rect -7440 1800 -7435 1820
rect -7465 1795 -7435 1800
rect -7285 1820 -7255 1825
rect -7285 1800 -7280 1820
rect -7260 1800 -7255 1820
rect -7285 1795 -7255 1800
rect -7460 1700 -7440 1795
rect -7280 1700 -7260 1795
rect -7465 1695 -7435 1700
rect -7465 1675 -7460 1695
rect -7440 1675 -7435 1695
rect -7465 1670 -7435 1675
rect -7285 1695 -7255 1700
rect -7285 1675 -7280 1695
rect -7260 1675 -7255 1695
rect -7285 1670 -7255 1675
rect -7460 1665 -7440 1670
rect -7280 1665 -7260 1670
rect -7600 1615 -7570 1620
rect -7600 1595 -7595 1615
rect -7575 1595 -7570 1615
rect -7600 1590 -7570 1595
rect -7595 1585 -7575 1590
rect -7235 1500 -7215 1845
rect -7100 1825 -7080 1830
rect -6920 1825 -6900 1830
rect -6740 1825 -6720 1830
rect -6560 1825 -6540 1830
rect -6380 1825 -6360 1830
rect -6200 1825 -6180 1830
rect -6020 1825 -6000 1830
rect -5840 1825 -5820 1830
rect -5660 1825 -5640 1830
rect -5480 1825 -5460 1830
rect -5300 1825 -5280 1830
rect -5120 1825 -5100 1830
rect -7105 1820 -7075 1825
rect -7105 1800 -7100 1820
rect -7080 1800 -7075 1820
rect -7105 1795 -7075 1800
rect -6925 1820 -6895 1825
rect -6925 1800 -6920 1820
rect -6900 1800 -6895 1820
rect -6925 1795 -6895 1800
rect -6745 1820 -6715 1825
rect -6745 1800 -6740 1820
rect -6720 1800 -6715 1820
rect -6745 1795 -6715 1800
rect -6565 1820 -6535 1825
rect -6565 1800 -6560 1820
rect -6540 1800 -6535 1820
rect -6565 1795 -6535 1800
rect -6385 1820 -6355 1825
rect -6385 1800 -6380 1820
rect -6360 1800 -6355 1820
rect -6385 1795 -6355 1800
rect -6205 1820 -6175 1825
rect -6205 1800 -6200 1820
rect -6180 1800 -6175 1820
rect -6205 1795 -6175 1800
rect -6025 1820 -5995 1825
rect -6025 1800 -6020 1820
rect -6000 1800 -5995 1820
rect -6025 1795 -5995 1800
rect -5845 1820 -5815 1825
rect -5845 1800 -5840 1820
rect -5820 1800 -5815 1820
rect -5845 1795 -5815 1800
rect -5665 1820 -5635 1825
rect -5665 1800 -5660 1820
rect -5640 1800 -5635 1820
rect -5665 1795 -5635 1800
rect -5485 1820 -5455 1825
rect -5485 1800 -5480 1820
rect -5460 1800 -5455 1820
rect -5485 1795 -5455 1800
rect -5305 1820 -5275 1825
rect -5305 1800 -5300 1820
rect -5280 1800 -5275 1820
rect -5305 1795 -5275 1800
rect -5125 1820 -5095 1825
rect -5125 1800 -5120 1820
rect -5100 1800 -5095 1820
rect -5125 1795 -5095 1800
rect -7100 1790 -7080 1795
rect -6920 1790 -6900 1795
rect -6740 1790 -6720 1795
rect -6560 1790 -6540 1795
rect -6380 1790 -6360 1795
rect -6200 1790 -6180 1795
rect -6020 1790 -6000 1795
rect -5840 1790 -5820 1795
rect -5660 1790 -5640 1795
rect -5480 1790 -5460 1795
rect -5300 1790 -5280 1795
rect -5120 1790 -5100 1795
rect -7145 1620 -7125 1625
rect -6965 1620 -6945 1625
rect -6785 1620 -6765 1625
rect -6605 1620 -6585 1625
rect -6425 1620 -6405 1625
rect -6245 1620 -6225 1625
rect -6065 1620 -6045 1625
rect -5885 1620 -5865 1625
rect -5705 1620 -5685 1625
rect -5525 1620 -5505 1625
rect -5345 1620 -5325 1625
rect -5165 1620 -5145 1625
rect -7150 1615 -7120 1620
rect -7150 1595 -7145 1615
rect -7125 1595 -7120 1615
rect -7150 1590 -7120 1595
rect -6970 1615 -6940 1620
rect -6970 1595 -6965 1615
rect -6945 1595 -6940 1615
rect -6970 1590 -6940 1595
rect -6790 1615 -6760 1620
rect -6790 1595 -6785 1615
rect -6765 1595 -6760 1615
rect -6790 1590 -6760 1595
rect -6610 1615 -6580 1620
rect -6610 1595 -6605 1615
rect -6585 1595 -6580 1615
rect -6610 1590 -6580 1595
rect -6430 1615 -6400 1620
rect -6430 1595 -6425 1615
rect -6405 1595 -6400 1615
rect -6430 1590 -6400 1595
rect -6250 1615 -6220 1620
rect -6250 1595 -6245 1615
rect -6225 1595 -6220 1615
rect -6250 1590 -6220 1595
rect -6070 1615 -6040 1620
rect -6070 1595 -6065 1615
rect -6045 1595 -6040 1615
rect -6070 1590 -6040 1595
rect -5890 1615 -5860 1620
rect -5890 1595 -5885 1615
rect -5865 1595 -5860 1615
rect -5890 1590 -5860 1595
rect -5710 1615 -5680 1620
rect -5710 1595 -5705 1615
rect -5685 1595 -5680 1615
rect -5710 1590 -5680 1595
rect -5530 1615 -5500 1620
rect -5530 1595 -5525 1615
rect -5505 1595 -5500 1615
rect -5530 1590 -5500 1595
rect -5350 1615 -5320 1620
rect -5350 1595 -5345 1615
rect -5325 1595 -5320 1615
rect -5350 1590 -5320 1595
rect -5170 1615 -5140 1620
rect -5170 1595 -5165 1615
rect -5145 1595 -5140 1615
rect -5170 1590 -5140 1595
rect -7190 1540 -7170 1545
rect -7195 1535 -7165 1540
rect -7195 1515 -7190 1535
rect -7170 1515 -7165 1535
rect -7195 1510 -7165 1515
rect -7240 1495 -7210 1500
rect -7240 1475 -7235 1495
rect -7215 1475 -7210 1495
rect -7240 1470 -7210 1475
rect -7235 1465 -7215 1470
rect -8270 1460 -8250 1465
rect -8090 1460 -8070 1465
rect -9715 1455 -9685 1460
rect -9715 1435 -9710 1455
rect -9690 1435 -9685 1455
rect -9715 1430 -9685 1435
rect -9535 1455 -9505 1460
rect -9535 1435 -9530 1455
rect -9510 1435 -9505 1455
rect -9535 1430 -9505 1435
rect -9355 1455 -9325 1460
rect -9355 1435 -9350 1455
rect -9330 1435 -9325 1455
rect -9355 1430 -9325 1435
rect -9175 1455 -9145 1460
rect -9175 1435 -9170 1455
rect -9150 1435 -9145 1455
rect -9175 1430 -9145 1435
rect -8680 1455 -8650 1460
rect -8680 1435 -8675 1455
rect -8655 1435 -8650 1455
rect -8680 1430 -8650 1435
rect -8275 1455 -8245 1460
rect -8275 1435 -8270 1455
rect -8250 1435 -8245 1455
rect -8275 1430 -8245 1435
rect -8095 1455 -8065 1460
rect -8095 1435 -8090 1455
rect -8070 1435 -8065 1455
rect -8095 1430 -8065 1435
rect -10070 1420 -10050 1425
rect -9890 1420 -9870 1425
rect -10075 1415 -10045 1420
rect -10075 1395 -10070 1415
rect -10050 1395 -10045 1415
rect -10075 1390 -10045 1395
rect -9895 1415 -9865 1420
rect -9895 1395 -9890 1415
rect -9870 1395 -9865 1415
rect -9895 1390 -9865 1395
rect -10070 1215 -10050 1390
rect -9890 1215 -9870 1390
rect -9710 1215 -9690 1430
rect -9530 1215 -9510 1430
rect -9350 1215 -9330 1430
rect -9170 1215 -9150 1430
rect -8990 1420 -8970 1425
rect -8810 1420 -8790 1425
rect -8995 1415 -8965 1420
rect -8995 1395 -8990 1415
rect -8970 1395 -8965 1415
rect -8995 1390 -8965 1395
rect -8815 1415 -8785 1420
rect -8815 1395 -8810 1415
rect -8790 1395 -8785 1415
rect -8815 1390 -8785 1395
rect -8990 1215 -8970 1390
rect -8810 1215 -8790 1390
rect -10075 1210 -10045 1215
rect -10075 1190 -10070 1210
rect -10050 1190 -10045 1210
rect -10075 1185 -10045 1190
rect -9895 1210 -9865 1215
rect -9895 1190 -9890 1210
rect -9870 1190 -9865 1210
rect -9895 1185 -9865 1190
rect -9715 1210 -9685 1215
rect -9715 1190 -9710 1210
rect -9690 1190 -9685 1210
rect -9715 1185 -9685 1190
rect -9535 1210 -9505 1215
rect -9535 1190 -9530 1210
rect -9510 1190 -9505 1210
rect -9535 1185 -9505 1190
rect -9355 1210 -9325 1215
rect -9355 1190 -9350 1210
rect -9330 1190 -9325 1210
rect -9355 1185 -9325 1190
rect -9175 1210 -9145 1215
rect -9175 1190 -9170 1210
rect -9150 1190 -9145 1210
rect -9175 1185 -9145 1190
rect -8995 1210 -8965 1215
rect -8995 1190 -8990 1210
rect -8970 1190 -8965 1210
rect -8995 1185 -8965 1190
rect -8815 1210 -8785 1215
rect -8815 1190 -8810 1210
rect -8790 1190 -8785 1210
rect -8815 1185 -8785 1190
rect -10070 1180 -10050 1185
rect -9890 1180 -9870 1185
rect -9710 1180 -9690 1185
rect -9530 1180 -9510 1185
rect -9350 1180 -9330 1185
rect -9170 1180 -9150 1185
rect -8990 1180 -8970 1185
rect -8810 1180 -8790 1185
rect -8675 1165 -8655 1430
rect -8630 1420 -8610 1425
rect -8450 1420 -8430 1425
rect -8635 1415 -8605 1420
rect -8635 1395 -8630 1415
rect -8610 1395 -8605 1415
rect -8635 1390 -8605 1395
rect -8455 1415 -8425 1420
rect -8455 1395 -8450 1415
rect -8430 1395 -8425 1415
rect -8455 1390 -8425 1395
rect -8630 1215 -8610 1390
rect -8450 1215 -8430 1390
rect -8270 1215 -8250 1430
rect -8090 1215 -8070 1430
rect -7550 1420 -7530 1425
rect -7370 1420 -7350 1425
rect -7555 1415 -7525 1420
rect -7555 1395 -7550 1415
rect -7530 1395 -7525 1415
rect -7555 1390 -7525 1395
rect -7375 1415 -7345 1420
rect -7375 1395 -7370 1415
rect -7350 1395 -7345 1415
rect -7375 1390 -7345 1395
rect -7910 1380 -7890 1385
rect -7730 1380 -7710 1385
rect -7915 1375 -7885 1380
rect -7915 1355 -7910 1375
rect -7890 1355 -7885 1375
rect -7915 1350 -7885 1355
rect -7735 1375 -7705 1380
rect -7735 1355 -7730 1375
rect -7710 1355 -7705 1375
rect -7735 1350 -7705 1355
rect -7910 1215 -7890 1350
rect -7730 1215 -7710 1350
rect -7550 1215 -7530 1390
rect -7370 1215 -7350 1390
rect -7235 1300 -7215 1305
rect -7240 1295 -7210 1300
rect -7240 1275 -7235 1295
rect -7215 1275 -7210 1295
rect -7240 1270 -7210 1275
rect -8635 1210 -8605 1215
rect -8635 1190 -8630 1210
rect -8610 1190 -8605 1210
rect -8635 1185 -8605 1190
rect -8455 1210 -8425 1215
rect -8455 1190 -8450 1210
rect -8430 1190 -8425 1210
rect -8455 1185 -8425 1190
rect -8275 1210 -8245 1215
rect -8275 1190 -8270 1210
rect -8250 1190 -8245 1210
rect -8275 1185 -8245 1190
rect -8095 1210 -8065 1215
rect -8095 1190 -8090 1210
rect -8070 1190 -8065 1210
rect -8095 1185 -8065 1190
rect -7915 1210 -7885 1215
rect -7915 1190 -7910 1210
rect -7890 1190 -7885 1210
rect -7915 1185 -7885 1190
rect -7735 1210 -7705 1215
rect -7735 1190 -7730 1210
rect -7710 1190 -7705 1210
rect -7735 1185 -7705 1190
rect -7555 1210 -7525 1215
rect -7555 1190 -7550 1210
rect -7530 1190 -7525 1210
rect -7555 1185 -7525 1190
rect -7375 1210 -7345 1215
rect -7375 1190 -7370 1210
rect -7350 1190 -7345 1210
rect -7375 1185 -7345 1190
rect -8630 1180 -8610 1185
rect -8450 1180 -8430 1185
rect -8270 1180 -8250 1185
rect -8090 1180 -8070 1185
rect -7910 1180 -7890 1185
rect -7730 1180 -7710 1185
rect -7550 1180 -7530 1185
rect -7370 1180 -7350 1185
rect -7235 1165 -7215 1270
rect -7190 1215 -7170 1510
rect -7195 1210 -7165 1215
rect -7195 1190 -7190 1210
rect -7170 1190 -7165 1210
rect -7195 1185 -7165 1190
rect -7190 1180 -7170 1185
rect -7145 1165 -7125 1590
rect -7010 1540 -6990 1545
rect -7015 1535 -6985 1540
rect -7015 1515 -7010 1535
rect -6990 1515 -6985 1535
rect -7015 1510 -6985 1515
rect -7055 1300 -7035 1305
rect -7060 1295 -7030 1300
rect -7060 1275 -7055 1295
rect -7035 1275 -7030 1295
rect -7060 1270 -7030 1275
rect -7055 1165 -7035 1270
rect -7010 1215 -6990 1510
rect -7015 1210 -6985 1215
rect -7015 1190 -7010 1210
rect -6990 1190 -6985 1210
rect -7015 1185 -6985 1190
rect -7010 1180 -6990 1185
rect -6965 1165 -6945 1590
rect -6830 1540 -6810 1545
rect -6835 1535 -6805 1540
rect -6835 1515 -6830 1535
rect -6810 1515 -6805 1535
rect -6835 1510 -6805 1515
rect -6875 1300 -6855 1305
rect -6880 1295 -6850 1300
rect -6880 1275 -6875 1295
rect -6855 1275 -6850 1295
rect -6880 1270 -6850 1275
rect -6875 1165 -6855 1270
rect -6830 1215 -6810 1510
rect -6835 1210 -6805 1215
rect -6835 1190 -6830 1210
rect -6810 1190 -6805 1210
rect -6835 1185 -6805 1190
rect -6830 1180 -6810 1185
rect -6785 1165 -6765 1590
rect -6650 1540 -6630 1545
rect -6655 1535 -6625 1540
rect -6655 1515 -6650 1535
rect -6630 1515 -6625 1535
rect -6655 1510 -6625 1515
rect -6695 1300 -6675 1305
rect -6700 1295 -6670 1300
rect -6700 1275 -6695 1295
rect -6675 1275 -6670 1295
rect -6700 1270 -6670 1275
rect -6695 1165 -6675 1270
rect -6650 1215 -6630 1510
rect -6655 1210 -6625 1215
rect -6655 1190 -6650 1210
rect -6630 1190 -6625 1210
rect -6655 1185 -6625 1190
rect -6650 1180 -6630 1185
rect -6605 1165 -6585 1590
rect -6470 1540 -6450 1545
rect -6475 1535 -6445 1540
rect -6475 1515 -6470 1535
rect -6450 1515 -6445 1535
rect -6475 1510 -6445 1515
rect -6515 1300 -6495 1305
rect -6520 1295 -6490 1300
rect -6520 1275 -6515 1295
rect -6495 1275 -6490 1295
rect -6520 1270 -6490 1275
rect -6515 1165 -6495 1270
rect -6470 1215 -6450 1510
rect -6475 1210 -6445 1215
rect -6475 1190 -6470 1210
rect -6450 1190 -6445 1210
rect -6475 1185 -6445 1190
rect -6470 1180 -6450 1185
rect -6425 1165 -6405 1590
rect -6290 1540 -6270 1545
rect -6295 1535 -6265 1540
rect -6295 1515 -6290 1535
rect -6270 1515 -6265 1535
rect -6295 1510 -6265 1515
rect -6335 1300 -6315 1305
rect -6340 1295 -6310 1300
rect -6340 1275 -6335 1295
rect -6315 1275 -6310 1295
rect -6340 1270 -6310 1275
rect -6335 1165 -6315 1270
rect -6290 1215 -6270 1510
rect -6295 1210 -6265 1215
rect -6295 1190 -6290 1210
rect -6270 1190 -6265 1210
rect -6295 1185 -6265 1190
rect -6290 1180 -6270 1185
rect -6245 1165 -6225 1590
rect -6110 1540 -6090 1545
rect -6115 1535 -6085 1540
rect -6115 1515 -6110 1535
rect -6090 1515 -6085 1535
rect -6115 1510 -6085 1515
rect -6155 1300 -6135 1305
rect -6160 1295 -6130 1300
rect -6160 1275 -6155 1295
rect -6135 1275 -6130 1295
rect -6160 1270 -6130 1275
rect -6155 1165 -6135 1270
rect -6110 1215 -6090 1510
rect -6115 1210 -6085 1215
rect -6115 1190 -6110 1210
rect -6090 1190 -6085 1210
rect -6115 1185 -6085 1190
rect -6110 1180 -6090 1185
rect -6065 1165 -6045 1590
rect -5930 1540 -5910 1545
rect -5935 1535 -5905 1540
rect -5935 1515 -5930 1535
rect -5910 1515 -5905 1535
rect -5935 1510 -5905 1515
rect -5975 1300 -5955 1305
rect -5980 1295 -5950 1300
rect -5980 1275 -5975 1295
rect -5955 1275 -5950 1295
rect -5980 1270 -5950 1275
rect -5975 1165 -5955 1270
rect -5930 1215 -5910 1510
rect -5935 1210 -5905 1215
rect -5935 1190 -5930 1210
rect -5910 1190 -5905 1210
rect -5935 1185 -5905 1190
rect -5930 1180 -5910 1185
rect -5885 1165 -5865 1590
rect -5750 1540 -5730 1545
rect -5755 1535 -5725 1540
rect -5755 1515 -5750 1535
rect -5730 1515 -5725 1535
rect -5755 1510 -5725 1515
rect -5795 1300 -5775 1305
rect -5800 1295 -5770 1300
rect -5800 1275 -5795 1295
rect -5775 1275 -5770 1295
rect -5800 1270 -5770 1275
rect -5795 1165 -5775 1270
rect -5750 1215 -5730 1510
rect -5755 1210 -5725 1215
rect -5755 1190 -5750 1210
rect -5730 1190 -5725 1210
rect -5755 1185 -5725 1190
rect -5750 1180 -5730 1185
rect -5705 1165 -5685 1590
rect -5570 1540 -5550 1545
rect -5575 1535 -5545 1540
rect -5575 1515 -5570 1535
rect -5550 1515 -5545 1535
rect -5575 1510 -5545 1515
rect -5615 1300 -5595 1305
rect -5620 1295 -5590 1300
rect -5620 1275 -5615 1295
rect -5595 1275 -5590 1295
rect -5620 1270 -5590 1275
rect -5615 1165 -5595 1270
rect -5570 1215 -5550 1510
rect -5575 1210 -5545 1215
rect -5575 1190 -5570 1210
rect -5550 1190 -5545 1210
rect -5575 1185 -5545 1190
rect -5570 1180 -5550 1185
rect -5525 1165 -5505 1590
rect -5390 1540 -5370 1545
rect -5395 1535 -5365 1540
rect -5395 1515 -5390 1535
rect -5370 1515 -5365 1535
rect -5395 1510 -5365 1515
rect -5435 1300 -5415 1305
rect -5440 1295 -5410 1300
rect -5440 1275 -5435 1295
rect -5415 1275 -5410 1295
rect -5440 1270 -5410 1275
rect -5435 1165 -5415 1270
rect -5390 1215 -5370 1510
rect -5395 1210 -5365 1215
rect -5395 1190 -5390 1210
rect -5370 1190 -5365 1210
rect -5395 1185 -5365 1190
rect -5390 1180 -5370 1185
rect -5345 1165 -5325 1590
rect -5210 1540 -5190 1545
rect -5215 1535 -5185 1540
rect -5215 1515 -5210 1535
rect -5190 1515 -5185 1535
rect -5215 1510 -5185 1515
rect -5255 1300 -5235 1305
rect -5260 1295 -5230 1300
rect -5260 1275 -5255 1295
rect -5235 1275 -5230 1295
rect -5260 1270 -5230 1275
rect -5255 1165 -5235 1270
rect -5210 1215 -5190 1510
rect -5215 1210 -5185 1215
rect -5215 1190 -5210 1210
rect -5190 1190 -5185 1210
rect -5215 1185 -5185 1190
rect -5210 1180 -5190 1185
rect -5165 1165 -5145 1590
rect -5075 1500 -5055 1845
rect -4940 1825 -4920 1830
rect -4760 1825 -4740 1830
rect -4945 1820 -4915 1825
rect -4945 1800 -4940 1820
rect -4920 1800 -4915 1820
rect -4945 1795 -4915 1800
rect -4765 1820 -4735 1825
rect -4765 1800 -4760 1820
rect -4740 1800 -4735 1820
rect -4765 1795 -4735 1800
rect -4940 1700 -4920 1795
rect -4760 1700 -4740 1795
rect -4945 1695 -4915 1700
rect -4945 1675 -4940 1695
rect -4920 1675 -4915 1695
rect -4945 1670 -4915 1675
rect -4765 1695 -4735 1700
rect -4765 1675 -4760 1695
rect -4740 1675 -4735 1695
rect -4765 1670 -4735 1675
rect -4940 1665 -4920 1670
rect -4760 1665 -4740 1670
rect -4715 1620 -4695 1845
rect -4580 1825 -4560 1830
rect -4400 1825 -4380 1830
rect -4220 1825 -4200 1830
rect -4040 1825 -4020 1830
rect -4585 1820 -4555 1825
rect -4585 1800 -4580 1820
rect -4560 1800 -4555 1820
rect -4585 1795 -4555 1800
rect -4405 1820 -4375 1825
rect -4405 1800 -4400 1820
rect -4380 1800 -4375 1820
rect -4405 1795 -4375 1800
rect -4225 1820 -4195 1825
rect -4225 1800 -4220 1820
rect -4200 1800 -4195 1820
rect -4225 1795 -4195 1800
rect -4045 1820 -4015 1825
rect -4045 1800 -4040 1820
rect -4020 1800 -4015 1820
rect -4045 1795 -4015 1800
rect -4580 1740 -4560 1795
rect -4400 1740 -4380 1795
rect -4220 1740 -4200 1795
rect -4040 1740 -4020 1795
rect -4585 1735 -4555 1740
rect -4585 1715 -4580 1735
rect -4560 1715 -4555 1735
rect -4585 1710 -4555 1715
rect -4405 1735 -4375 1740
rect -4405 1715 -4400 1735
rect -4380 1715 -4375 1735
rect -4405 1710 -4375 1715
rect -4225 1735 -4195 1740
rect -4225 1715 -4220 1735
rect -4200 1715 -4195 1735
rect -4225 1710 -4195 1715
rect -4045 1735 -4015 1740
rect -4045 1715 -4040 1735
rect -4020 1715 -4015 1735
rect -4045 1710 -4015 1715
rect -4580 1705 -4560 1710
rect -4400 1705 -4380 1710
rect -4220 1705 -4200 1710
rect -4040 1705 -4020 1710
rect -3995 1660 -3975 1845
rect -3860 1825 -3840 1830
rect -3680 1825 -3660 1830
rect -3865 1820 -3835 1825
rect -3865 1800 -3860 1820
rect -3840 1800 -3835 1820
rect -3865 1795 -3835 1800
rect -3685 1820 -3655 1825
rect -3685 1800 -3680 1820
rect -3660 1800 -3655 1820
rect -3685 1795 -3655 1800
rect -3860 1700 -3840 1795
rect -3680 1700 -3660 1795
rect -3865 1695 -3835 1700
rect -3865 1675 -3860 1695
rect -3840 1675 -3835 1695
rect -3865 1670 -3835 1675
rect -3685 1695 -3655 1700
rect -3685 1675 -3680 1695
rect -3660 1675 -3655 1695
rect -3685 1670 -3655 1675
rect -3860 1665 -3840 1670
rect -3680 1665 -3660 1670
rect -4000 1655 -3970 1660
rect -4000 1635 -3995 1655
rect -3975 1635 -3970 1655
rect -4000 1630 -3970 1635
rect -3995 1625 -3975 1630
rect -4720 1615 -4690 1620
rect -4720 1595 -4715 1615
rect -4695 1595 -4690 1615
rect -4720 1590 -4690 1595
rect -4715 1585 -4695 1590
rect -5080 1495 -5050 1500
rect -5080 1475 -5075 1495
rect -5055 1475 -5050 1495
rect -5080 1470 -5050 1475
rect -5075 1465 -5055 1470
rect -3635 1460 -3615 1845
rect -3500 1825 -3480 1830
rect -3320 1825 -3300 1830
rect -3140 1825 -3120 1830
rect -2960 1825 -2940 1830
rect -2780 1825 -2760 1830
rect -2600 1825 -2580 1830
rect -2420 1825 -2400 1830
rect -2240 1825 -2220 1830
rect -2060 1825 -2040 1830
rect -1880 1825 -1860 1830
rect -1700 1825 -1680 1830
rect -1520 1825 -1500 1830
rect -3505 1820 -3475 1825
rect -3505 1800 -3500 1820
rect -3480 1800 -3475 1820
rect -3505 1795 -3475 1800
rect -3325 1820 -3295 1825
rect -3325 1800 -3320 1820
rect -3300 1800 -3295 1820
rect -3325 1795 -3295 1800
rect -3145 1820 -3115 1825
rect -3145 1800 -3140 1820
rect -3120 1800 -3115 1820
rect -3145 1795 -3115 1800
rect -2965 1820 -2935 1825
rect -2965 1800 -2960 1820
rect -2940 1800 -2935 1820
rect -2965 1795 -2935 1800
rect -2785 1820 -2755 1825
rect -2785 1800 -2780 1820
rect -2760 1800 -2755 1820
rect -2785 1795 -2755 1800
rect -2605 1820 -2575 1825
rect -2605 1800 -2600 1820
rect -2580 1800 -2575 1820
rect -2605 1795 -2575 1800
rect -2425 1820 -2395 1825
rect -2425 1800 -2420 1820
rect -2400 1800 -2395 1820
rect -2425 1795 -2395 1800
rect -2245 1820 -2215 1825
rect -2245 1800 -2240 1820
rect -2220 1800 -2215 1820
rect -2245 1795 -2215 1800
rect -2065 1820 -2035 1825
rect -2065 1800 -2060 1820
rect -2040 1800 -2035 1820
rect -2065 1795 -2035 1800
rect -1885 1820 -1855 1825
rect -1885 1800 -1880 1820
rect -1860 1800 -1855 1820
rect -1885 1795 -1855 1800
rect -1705 1820 -1675 1825
rect -1705 1800 -1700 1820
rect -1680 1800 -1675 1820
rect -1705 1795 -1675 1800
rect -1525 1820 -1495 1825
rect -1525 1800 -1520 1820
rect -1500 1800 -1495 1820
rect -1525 1795 -1495 1800
rect -3500 1790 -3480 1795
rect -3320 1790 -3300 1795
rect -3140 1790 -3120 1795
rect -2960 1790 -2940 1795
rect -2780 1790 -2760 1795
rect -2600 1790 -2580 1795
rect -2420 1790 -2400 1795
rect -2240 1790 -2220 1795
rect -2060 1790 -2040 1795
rect -1880 1790 -1860 1795
rect -1700 1790 -1680 1795
rect -1520 1790 -1500 1795
rect -3545 1660 -3525 1665
rect -3365 1660 -3345 1665
rect -3185 1660 -3165 1665
rect -3005 1660 -2985 1665
rect -2825 1660 -2805 1665
rect -2645 1660 -2625 1665
rect -2465 1660 -2445 1665
rect -2285 1660 -2265 1665
rect -2105 1660 -2085 1665
rect -1925 1660 -1905 1665
rect -1745 1660 -1725 1665
rect -1565 1660 -1545 1665
rect -3550 1655 -3520 1660
rect -3550 1635 -3545 1655
rect -3525 1635 -3520 1655
rect -3550 1630 -3520 1635
rect -3370 1655 -3340 1660
rect -3370 1635 -3365 1655
rect -3345 1635 -3340 1655
rect -3370 1630 -3340 1635
rect -3190 1655 -3160 1660
rect -3190 1635 -3185 1655
rect -3165 1635 -3160 1655
rect -3190 1630 -3160 1635
rect -3010 1655 -2980 1660
rect -3010 1635 -3005 1655
rect -2985 1635 -2980 1655
rect -3010 1630 -2980 1635
rect -2830 1655 -2800 1660
rect -2830 1635 -2825 1655
rect -2805 1635 -2800 1655
rect -2830 1630 -2800 1635
rect -2650 1655 -2620 1660
rect -2650 1635 -2645 1655
rect -2625 1635 -2620 1655
rect -2650 1630 -2620 1635
rect -2470 1655 -2440 1660
rect -2470 1635 -2465 1655
rect -2445 1635 -2440 1655
rect -2470 1630 -2440 1635
rect -2290 1655 -2260 1660
rect -2290 1635 -2285 1655
rect -2265 1635 -2260 1655
rect -2290 1630 -2260 1635
rect -2110 1655 -2080 1660
rect -2110 1635 -2105 1655
rect -2085 1635 -2080 1655
rect -2110 1630 -2080 1635
rect -1930 1655 -1900 1660
rect -1930 1635 -1925 1655
rect -1905 1635 -1900 1655
rect -1930 1630 -1900 1635
rect -1750 1655 -1720 1660
rect -1750 1635 -1745 1655
rect -1725 1635 -1720 1655
rect -1750 1630 -1720 1635
rect -1570 1655 -1540 1660
rect -1570 1635 -1565 1655
rect -1545 1635 -1540 1655
rect -1570 1630 -1540 1635
rect -3590 1580 -3570 1585
rect -3595 1575 -3565 1580
rect -3595 1555 -3590 1575
rect -3570 1555 -3565 1575
rect -3595 1550 -3565 1555
rect -3640 1455 -3610 1460
rect -3640 1435 -3635 1455
rect -3615 1435 -3610 1455
rect -3640 1430 -3610 1435
rect -3635 1425 -3615 1430
rect -5030 1420 -5010 1425
rect -4850 1420 -4830 1425
rect -3950 1420 -3930 1425
rect -3770 1420 -3750 1425
rect -5035 1415 -5005 1420
rect -5035 1395 -5030 1415
rect -5010 1395 -5005 1415
rect -5035 1390 -5005 1395
rect -4855 1415 -4825 1420
rect -4855 1395 -4850 1415
rect -4830 1395 -4825 1415
rect -4855 1390 -4825 1395
rect -3955 1415 -3925 1420
rect -3955 1395 -3950 1415
rect -3930 1395 -3925 1415
rect -3955 1390 -3925 1395
rect -3775 1415 -3745 1420
rect -3775 1395 -3770 1415
rect -3750 1395 -3745 1415
rect -3775 1390 -3745 1395
rect -5075 1300 -5055 1305
rect -5080 1295 -5050 1300
rect -5080 1275 -5075 1295
rect -5055 1275 -5050 1295
rect -5080 1270 -5050 1275
rect -5075 1165 -5055 1270
rect -5030 1215 -5010 1390
rect -4850 1215 -4830 1390
rect -4670 1380 -4650 1385
rect -4490 1380 -4470 1385
rect -4310 1380 -4290 1385
rect -4130 1380 -4110 1385
rect -4675 1375 -4645 1380
rect -4675 1355 -4670 1375
rect -4650 1355 -4645 1375
rect -4675 1350 -4645 1355
rect -4495 1375 -4465 1380
rect -4495 1355 -4490 1375
rect -4470 1355 -4465 1375
rect -4495 1350 -4465 1355
rect -4315 1375 -4285 1380
rect -4315 1355 -4310 1375
rect -4290 1355 -4285 1375
rect -4315 1350 -4285 1355
rect -4135 1375 -4105 1380
rect -4135 1355 -4130 1375
rect -4110 1355 -4105 1375
rect -4135 1350 -4105 1355
rect -4670 1215 -4650 1350
rect -4490 1215 -4470 1350
rect -4310 1215 -4290 1350
rect -4130 1215 -4110 1350
rect -3950 1215 -3930 1390
rect -3770 1215 -3750 1390
rect -3635 1300 -3615 1305
rect -3640 1295 -3610 1300
rect -3640 1275 -3635 1295
rect -3615 1275 -3610 1295
rect -3640 1270 -3610 1275
rect -5035 1210 -5005 1215
rect -5035 1190 -5030 1210
rect -5010 1190 -5005 1210
rect -5035 1185 -5005 1190
rect -4855 1210 -4825 1215
rect -4855 1190 -4850 1210
rect -4830 1190 -4825 1210
rect -4855 1185 -4825 1190
rect -4675 1210 -4645 1215
rect -4675 1190 -4670 1210
rect -4650 1190 -4645 1210
rect -4675 1185 -4645 1190
rect -4495 1210 -4465 1215
rect -4495 1190 -4490 1210
rect -4470 1190 -4465 1210
rect -4495 1185 -4465 1190
rect -4315 1210 -4285 1215
rect -4315 1190 -4310 1210
rect -4290 1190 -4285 1210
rect -4315 1185 -4285 1190
rect -4135 1210 -4105 1215
rect -4135 1190 -4130 1210
rect -4110 1190 -4105 1210
rect -4135 1185 -4105 1190
rect -3955 1210 -3925 1215
rect -3955 1190 -3950 1210
rect -3930 1190 -3925 1210
rect -3955 1185 -3925 1190
rect -3775 1210 -3745 1215
rect -3775 1190 -3770 1210
rect -3750 1190 -3745 1210
rect -3775 1185 -3745 1190
rect -5030 1180 -5010 1185
rect -4850 1180 -4830 1185
rect -4670 1180 -4650 1185
rect -4490 1180 -4470 1185
rect -4310 1180 -4290 1185
rect -4130 1180 -4110 1185
rect -3950 1180 -3930 1185
rect -3770 1180 -3750 1185
rect -3635 1165 -3615 1270
rect -3590 1215 -3570 1550
rect -3595 1210 -3565 1215
rect -3595 1190 -3590 1210
rect -3570 1190 -3565 1210
rect -3595 1185 -3565 1190
rect -3590 1180 -3570 1185
rect -3545 1165 -3525 1630
rect -3410 1580 -3390 1585
rect -3415 1575 -3385 1580
rect -3415 1555 -3410 1575
rect -3390 1555 -3385 1575
rect -3415 1550 -3385 1555
rect -3455 1300 -3435 1305
rect -3460 1295 -3430 1300
rect -3460 1275 -3455 1295
rect -3435 1275 -3430 1295
rect -3460 1270 -3430 1275
rect -3455 1165 -3435 1270
rect -3410 1215 -3390 1550
rect -3415 1210 -3385 1215
rect -3415 1190 -3410 1210
rect -3390 1190 -3385 1210
rect -3415 1185 -3385 1190
rect -3410 1180 -3390 1185
rect -3365 1165 -3345 1630
rect -3230 1580 -3210 1585
rect -3235 1575 -3205 1580
rect -3235 1555 -3230 1575
rect -3210 1555 -3205 1575
rect -3235 1550 -3205 1555
rect -3275 1300 -3255 1305
rect -3280 1295 -3250 1300
rect -3280 1275 -3275 1295
rect -3255 1275 -3250 1295
rect -3280 1270 -3250 1275
rect -3275 1165 -3255 1270
rect -3230 1215 -3210 1550
rect -3235 1210 -3205 1215
rect -3235 1190 -3230 1210
rect -3210 1190 -3205 1210
rect -3235 1185 -3205 1190
rect -3230 1180 -3210 1185
rect -3185 1165 -3165 1630
rect -3050 1580 -3030 1585
rect -3055 1575 -3025 1580
rect -3055 1555 -3050 1575
rect -3030 1555 -3025 1575
rect -3055 1550 -3025 1555
rect -3095 1300 -3075 1305
rect -3100 1295 -3070 1300
rect -3100 1275 -3095 1295
rect -3075 1275 -3070 1295
rect -3100 1270 -3070 1275
rect -3095 1165 -3075 1270
rect -3050 1215 -3030 1550
rect -3055 1210 -3025 1215
rect -3055 1190 -3050 1210
rect -3030 1190 -3025 1210
rect -3055 1185 -3025 1190
rect -3050 1180 -3030 1185
rect -3005 1165 -2985 1630
rect -2870 1580 -2850 1585
rect -2875 1575 -2845 1580
rect -2875 1555 -2870 1575
rect -2850 1555 -2845 1575
rect -2875 1550 -2845 1555
rect -2915 1300 -2895 1305
rect -2920 1295 -2890 1300
rect -2920 1275 -2915 1295
rect -2895 1275 -2890 1295
rect -2920 1270 -2890 1275
rect -2915 1165 -2895 1270
rect -2870 1215 -2850 1550
rect -2875 1210 -2845 1215
rect -2875 1190 -2870 1210
rect -2850 1190 -2845 1210
rect -2875 1185 -2845 1190
rect -2870 1180 -2850 1185
rect -2825 1165 -2805 1630
rect -2690 1580 -2670 1585
rect -2695 1575 -2665 1580
rect -2695 1555 -2690 1575
rect -2670 1555 -2665 1575
rect -2695 1550 -2665 1555
rect -2735 1300 -2715 1305
rect -2740 1295 -2710 1300
rect -2740 1275 -2735 1295
rect -2715 1275 -2710 1295
rect -2740 1270 -2710 1275
rect -2735 1165 -2715 1270
rect -2690 1215 -2670 1550
rect -2695 1210 -2665 1215
rect -2695 1190 -2690 1210
rect -2670 1190 -2665 1210
rect -2695 1185 -2665 1190
rect -2690 1180 -2670 1185
rect -2645 1165 -2625 1630
rect -2510 1580 -2490 1585
rect -2515 1575 -2485 1580
rect -2515 1555 -2510 1575
rect -2490 1555 -2485 1575
rect -2515 1550 -2485 1555
rect -2555 1300 -2535 1305
rect -2560 1295 -2530 1300
rect -2560 1275 -2555 1295
rect -2535 1275 -2530 1295
rect -2560 1270 -2530 1275
rect -2555 1165 -2535 1270
rect -2510 1215 -2490 1550
rect -2515 1210 -2485 1215
rect -2515 1190 -2510 1210
rect -2490 1190 -2485 1210
rect -2515 1185 -2485 1190
rect -2510 1180 -2490 1185
rect -2465 1165 -2445 1630
rect -2330 1580 -2310 1585
rect -2335 1575 -2305 1580
rect -2335 1555 -2330 1575
rect -2310 1555 -2305 1575
rect -2335 1550 -2305 1555
rect -2375 1300 -2355 1305
rect -2380 1295 -2350 1300
rect -2380 1275 -2375 1295
rect -2355 1275 -2350 1295
rect -2380 1270 -2350 1275
rect -2375 1165 -2355 1270
rect -2330 1215 -2310 1550
rect -2335 1210 -2305 1215
rect -2335 1190 -2330 1210
rect -2310 1190 -2305 1210
rect -2335 1185 -2305 1190
rect -2330 1180 -2310 1185
rect -2285 1165 -2265 1630
rect -2150 1580 -2130 1585
rect -2155 1575 -2125 1580
rect -2155 1555 -2150 1575
rect -2130 1555 -2125 1575
rect -2155 1550 -2125 1555
rect -2195 1300 -2175 1305
rect -2200 1295 -2170 1300
rect -2200 1275 -2195 1295
rect -2175 1275 -2170 1295
rect -2200 1270 -2170 1275
rect -2195 1165 -2175 1270
rect -2150 1215 -2130 1550
rect -2155 1210 -2125 1215
rect -2155 1190 -2150 1210
rect -2130 1190 -2125 1210
rect -2155 1185 -2125 1190
rect -2150 1180 -2130 1185
rect -2105 1165 -2085 1630
rect -1970 1580 -1950 1585
rect -1975 1575 -1945 1580
rect -1975 1555 -1970 1575
rect -1950 1555 -1945 1575
rect -1975 1550 -1945 1555
rect -2015 1300 -1995 1305
rect -2020 1295 -1990 1300
rect -2020 1275 -2015 1295
rect -1995 1275 -1990 1295
rect -2020 1270 -1990 1275
rect -2015 1165 -1995 1270
rect -1970 1215 -1950 1550
rect -1975 1210 -1945 1215
rect -1975 1190 -1970 1210
rect -1950 1190 -1945 1210
rect -1975 1185 -1945 1190
rect -1970 1180 -1950 1185
rect -1925 1165 -1905 1630
rect -1790 1580 -1770 1585
rect -1795 1575 -1765 1580
rect -1795 1555 -1790 1575
rect -1770 1555 -1765 1575
rect -1795 1550 -1765 1555
rect -1835 1300 -1815 1305
rect -1840 1295 -1810 1300
rect -1840 1275 -1835 1295
rect -1815 1275 -1810 1295
rect -1840 1270 -1810 1275
rect -1835 1165 -1815 1270
rect -1790 1215 -1770 1550
rect -1795 1210 -1765 1215
rect -1795 1190 -1790 1210
rect -1770 1190 -1765 1210
rect -1795 1185 -1765 1190
rect -1790 1180 -1770 1185
rect -1745 1165 -1725 1630
rect -1610 1580 -1590 1585
rect -1615 1575 -1585 1580
rect -1615 1555 -1610 1575
rect -1590 1555 -1585 1575
rect -1615 1550 -1585 1555
rect -1655 1300 -1635 1305
rect -1660 1295 -1630 1300
rect -1660 1275 -1655 1295
rect -1635 1275 -1630 1295
rect -1660 1270 -1630 1275
rect -1655 1165 -1635 1270
rect -1610 1215 -1590 1550
rect -1615 1210 -1585 1215
rect -1615 1190 -1610 1210
rect -1590 1190 -1585 1210
rect -1615 1185 -1585 1190
rect -1610 1180 -1590 1185
rect -1565 1165 -1545 1630
rect -1475 1460 -1455 1845
rect -1340 1825 -1320 1830
rect -1160 1825 -1140 1830
rect -1345 1820 -1315 1825
rect -1345 1800 -1340 1820
rect -1320 1800 -1315 1820
rect -1345 1795 -1315 1800
rect -1165 1820 -1135 1825
rect -1165 1800 -1160 1820
rect -1140 1800 -1135 1820
rect -1165 1795 -1135 1800
rect -1340 1700 -1320 1795
rect -1160 1700 -1140 1795
rect -1345 1695 -1315 1700
rect -1345 1675 -1340 1695
rect -1320 1675 -1315 1695
rect -1345 1670 -1315 1675
rect -1165 1695 -1135 1700
rect -1165 1675 -1160 1695
rect -1140 1675 -1135 1695
rect -1165 1670 -1135 1675
rect -1340 1665 -1320 1670
rect -1160 1665 -1140 1670
rect -1115 1660 -1095 1845
rect -980 1825 -960 1830
rect -800 1825 -780 1830
rect -985 1820 -955 1825
rect -985 1800 -980 1820
rect -960 1800 -955 1820
rect -985 1795 -955 1800
rect -805 1820 -775 1825
rect -805 1800 -800 1820
rect -780 1800 -775 1820
rect -805 1795 -775 1800
rect -980 1740 -960 1795
rect -800 1740 -780 1795
rect -985 1735 -955 1740
rect -985 1715 -980 1735
rect -960 1715 -955 1735
rect -985 1710 -955 1715
rect -805 1735 -775 1740
rect -805 1715 -800 1735
rect -780 1715 -775 1735
rect -805 1710 -775 1715
rect -980 1705 -960 1710
rect -800 1705 -780 1710
rect -1120 1655 -1090 1660
rect -1120 1635 -1115 1655
rect -1095 1635 -1090 1655
rect -1120 1630 -1090 1635
rect -1115 1625 -1095 1630
rect -1480 1455 -1450 1460
rect -1480 1435 -1475 1455
rect -1455 1435 -1450 1455
rect -1480 1430 -1450 1435
rect -1475 1425 -1455 1430
rect -1430 1420 -1410 1425
rect -1250 1420 -1230 1425
rect -1435 1415 -1405 1420
rect -1435 1395 -1430 1415
rect -1410 1395 -1405 1415
rect -1435 1390 -1405 1395
rect -1255 1415 -1225 1420
rect -1255 1395 -1250 1415
rect -1230 1395 -1225 1415
rect -1255 1390 -1225 1395
rect -1475 1300 -1455 1305
rect -1480 1295 -1450 1300
rect -1480 1275 -1475 1295
rect -1455 1275 -1450 1295
rect -1480 1270 -1450 1275
rect -1475 1165 -1455 1270
rect -1430 1215 -1410 1390
rect -1250 1215 -1230 1390
rect -1070 1380 -1050 1385
rect -890 1380 -870 1385
rect -1075 1375 -1045 1380
rect -1075 1355 -1070 1375
rect -1050 1355 -1045 1375
rect -1075 1350 -1045 1355
rect -895 1375 -865 1380
rect -895 1355 -890 1375
rect -870 1355 -865 1375
rect -895 1350 -865 1355
rect -1070 1215 -1050 1350
rect -890 1215 -870 1350
rect -1435 1210 -1405 1215
rect -1435 1190 -1430 1210
rect -1410 1190 -1405 1210
rect -1435 1185 -1405 1190
rect -1255 1210 -1225 1215
rect -1255 1190 -1250 1210
rect -1230 1190 -1225 1210
rect -1255 1185 -1225 1190
rect -1075 1210 -1045 1215
rect -1075 1190 -1070 1210
rect -1050 1190 -1045 1210
rect -1075 1185 -1045 1190
rect -895 1210 -865 1215
rect -895 1190 -890 1210
rect -870 1190 -865 1210
rect -895 1185 -865 1190
rect -1430 1180 -1410 1185
rect -1250 1180 -1230 1185
rect -1070 1180 -1050 1185
rect -890 1180 -870 1185
rect -665 1165 -645 1845
rect -575 1300 -555 1845
rect -485 1460 -465 1845
rect -490 1455 -460 1460
rect -490 1435 -485 1455
rect -465 1435 -460 1455
rect -490 1430 -460 1435
rect -580 1295 -550 1300
rect -580 1275 -575 1295
rect -555 1275 -550 1295
rect -580 1270 -550 1275
rect -575 1165 -555 1270
rect -485 1165 -465 1430
rect -395 1380 -375 1845
rect -305 1420 -285 1845
rect -215 1700 -195 1845
rect -125 1740 -105 1845
rect -130 1735 -100 1740
rect -130 1715 -125 1735
rect -105 1715 -100 1735
rect -130 1710 -100 1715
rect -220 1695 -190 1700
rect -220 1675 -215 1695
rect -195 1675 -190 1695
rect -220 1670 -190 1675
rect -310 1415 -280 1420
rect -310 1395 -305 1415
rect -285 1395 -280 1415
rect -310 1390 -280 1395
rect -400 1375 -370 1380
rect -400 1355 -395 1375
rect -375 1355 -370 1375
rect -400 1350 -370 1355
rect -395 1165 -375 1350
rect -305 1165 -285 1390
rect -215 1165 -195 1670
rect -125 1165 -105 1710
rect -11560 1155 -11530 1165
rect -11560 1075 -11555 1155
rect -11535 1075 -11530 1155
rect -11560 1065 -11530 1075
rect -11470 1065 -11440 1165
rect -11380 1065 -11350 1165
rect -11290 1065 -11260 1165
rect -11200 1065 -11170 1165
rect -11110 1065 -11080 1165
rect -11020 1065 -10990 1165
rect -10930 1065 -10900 1165
rect -10840 1155 -10810 1165
rect -10840 1075 -10835 1155
rect -10815 1075 -10810 1155
rect -10840 1065 -10810 1075
rect -10750 1155 -10720 1165
rect -10750 1075 -10745 1155
rect -10725 1075 -10720 1155
rect -10750 1065 -10720 1075
rect -10660 1155 -10630 1165
rect -10660 1075 -10655 1155
rect -10635 1075 -10630 1155
rect -10660 1065 -10630 1075
rect -10570 1155 -10540 1165
rect -10570 1075 -10565 1155
rect -10545 1075 -10540 1155
rect -10570 1065 -10540 1075
rect -10480 1155 -10450 1165
rect -10480 1075 -10475 1155
rect -10455 1075 -10450 1155
rect -10480 1065 -10450 1075
rect -10390 1155 -10360 1165
rect -10390 1075 -10385 1155
rect -10365 1075 -10360 1155
rect -10390 1065 -10360 1075
rect -10300 1155 -10270 1165
rect -10300 1075 -10295 1155
rect -10275 1075 -10270 1155
rect -10300 1065 -10270 1075
rect -10210 1155 -10180 1165
rect -10210 1075 -10205 1155
rect -10185 1075 -10180 1155
rect -10210 1065 -10180 1075
rect -10120 1155 -10090 1165
rect -10120 1075 -10115 1155
rect -10095 1075 -10090 1155
rect -10120 1065 -10090 1075
rect -10030 1155 -10000 1165
rect -10030 1075 -10025 1155
rect -10005 1075 -10000 1155
rect -10030 1065 -10000 1075
rect -9940 1155 -9910 1165
rect -9940 1075 -9935 1155
rect -9915 1075 -9910 1155
rect -9940 1065 -9910 1075
rect -9850 1155 -9820 1165
rect -9850 1075 -9845 1155
rect -9825 1075 -9820 1155
rect -9850 1065 -9820 1075
rect -9760 1155 -9730 1165
rect -9760 1075 -9755 1155
rect -9735 1075 -9730 1155
rect -9760 1065 -9730 1075
rect -9670 1155 -9640 1165
rect -9670 1075 -9665 1155
rect -9645 1075 -9640 1155
rect -9670 1065 -9640 1075
rect -9580 1155 -9550 1165
rect -9580 1075 -9575 1155
rect -9555 1075 -9550 1155
rect -9580 1065 -9550 1075
rect -9490 1155 -9460 1165
rect -9490 1075 -9485 1155
rect -9465 1075 -9460 1155
rect -9490 1065 -9460 1075
rect -9400 1155 -9370 1165
rect -9400 1075 -9395 1155
rect -9375 1075 -9370 1155
rect -9400 1065 -9370 1075
rect -9310 1155 -9280 1165
rect -9310 1075 -9305 1155
rect -9285 1075 -9280 1155
rect -9310 1065 -9280 1075
rect -9220 1155 -9190 1165
rect -9220 1075 -9215 1155
rect -9195 1075 -9190 1155
rect -9220 1065 -9190 1075
rect -9130 1155 -9100 1165
rect -9130 1075 -9125 1155
rect -9105 1075 -9100 1155
rect -9130 1065 -9100 1075
rect -9040 1155 -9010 1165
rect -9040 1075 -9035 1155
rect -9015 1075 -9010 1155
rect -9040 1065 -9010 1075
rect -8950 1155 -8920 1165
rect -8950 1075 -8945 1155
rect -8925 1075 -8920 1155
rect -8950 1065 -8920 1075
rect -8860 1155 -8830 1165
rect -8860 1075 -8855 1155
rect -8835 1075 -8830 1155
rect -8860 1065 -8830 1075
rect -8770 1155 -8740 1165
rect -8770 1075 -8765 1155
rect -8745 1075 -8740 1155
rect -8770 1065 -8740 1075
rect -8680 1155 -8650 1165
rect -8680 1075 -8675 1155
rect -8655 1075 -8650 1155
rect -8680 1065 -8650 1075
rect -8590 1155 -8560 1165
rect -8590 1075 -8585 1155
rect -8565 1075 -8560 1155
rect -8590 1065 -8560 1075
rect -8500 1155 -8470 1165
rect -8500 1075 -8495 1155
rect -8475 1075 -8470 1155
rect -8500 1065 -8470 1075
rect -8410 1155 -8380 1165
rect -8410 1075 -8405 1155
rect -8385 1075 -8380 1155
rect -8410 1065 -8380 1075
rect -8320 1155 -8290 1165
rect -8320 1075 -8315 1155
rect -8295 1075 -8290 1155
rect -8320 1065 -8290 1075
rect -8230 1155 -8200 1165
rect -8230 1075 -8225 1155
rect -8205 1075 -8200 1155
rect -8230 1065 -8200 1075
rect -8140 1155 -8110 1165
rect -8140 1075 -8135 1155
rect -8115 1075 -8110 1155
rect -8140 1065 -8110 1075
rect -8050 1155 -8020 1165
rect -8050 1075 -8045 1155
rect -8025 1075 -8020 1155
rect -8050 1065 -8020 1075
rect -7960 1155 -7930 1165
rect -7960 1075 -7955 1155
rect -7935 1075 -7930 1155
rect -7960 1065 -7930 1075
rect -7870 1155 -7840 1165
rect -7870 1075 -7865 1155
rect -7845 1075 -7840 1155
rect -7870 1065 -7840 1075
rect -7780 1155 -7750 1165
rect -7780 1075 -7775 1155
rect -7755 1075 -7750 1155
rect -7780 1065 -7750 1075
rect -7690 1155 -7660 1165
rect -7690 1075 -7685 1155
rect -7665 1075 -7660 1155
rect -7690 1065 -7660 1075
rect -7600 1155 -7570 1165
rect -7600 1075 -7595 1155
rect -7575 1075 -7570 1155
rect -7600 1065 -7570 1075
rect -7510 1155 -7480 1165
rect -7510 1075 -7505 1155
rect -7485 1075 -7480 1155
rect -7510 1065 -7480 1075
rect -7420 1155 -7390 1165
rect -7420 1075 -7415 1155
rect -7395 1075 -7390 1155
rect -7420 1065 -7390 1075
rect -7330 1155 -7300 1165
rect -7330 1075 -7325 1155
rect -7305 1075 -7300 1155
rect -7330 1065 -7300 1075
rect -7240 1155 -7210 1165
rect -7240 1075 -7235 1155
rect -7215 1075 -7210 1155
rect -7240 1065 -7210 1075
rect -7150 1155 -7120 1165
rect -7150 1075 -7145 1155
rect -7125 1075 -7120 1155
rect -7150 1065 -7120 1075
rect -7060 1155 -7030 1165
rect -7060 1075 -7055 1155
rect -7035 1075 -7030 1155
rect -7060 1065 -7030 1075
rect -6970 1155 -6940 1165
rect -6970 1075 -6965 1155
rect -6945 1075 -6940 1155
rect -6970 1065 -6940 1075
rect -6880 1155 -6850 1165
rect -6880 1075 -6875 1155
rect -6855 1075 -6850 1155
rect -6880 1065 -6850 1075
rect -6790 1155 -6760 1165
rect -6790 1075 -6785 1155
rect -6765 1075 -6760 1155
rect -6790 1065 -6760 1075
rect -6700 1155 -6670 1165
rect -6700 1075 -6695 1155
rect -6675 1075 -6670 1155
rect -6700 1065 -6670 1075
rect -6610 1155 -6580 1165
rect -6610 1075 -6605 1155
rect -6585 1075 -6580 1155
rect -6610 1065 -6580 1075
rect -6520 1155 -6490 1165
rect -6520 1075 -6515 1155
rect -6495 1075 -6490 1155
rect -6520 1065 -6490 1075
rect -6430 1155 -6400 1165
rect -6430 1075 -6425 1155
rect -6405 1075 -6400 1155
rect -6430 1065 -6400 1075
rect -6340 1155 -6310 1165
rect -6340 1075 -6335 1155
rect -6315 1075 -6310 1155
rect -6340 1065 -6310 1075
rect -6250 1155 -6220 1165
rect -6250 1075 -6245 1155
rect -6225 1075 -6220 1155
rect -6250 1065 -6220 1075
rect -6160 1155 -6130 1165
rect -6160 1075 -6155 1155
rect -6135 1075 -6130 1155
rect -6160 1065 -6130 1075
rect -6070 1155 -6040 1165
rect -6070 1075 -6065 1155
rect -6045 1075 -6040 1155
rect -6070 1065 -6040 1075
rect -5980 1155 -5950 1165
rect -5980 1075 -5975 1155
rect -5955 1075 -5950 1155
rect -5980 1065 -5950 1075
rect -5890 1155 -5860 1165
rect -5890 1075 -5885 1155
rect -5865 1075 -5860 1155
rect -5890 1065 -5860 1075
rect -5800 1155 -5770 1165
rect -5800 1075 -5795 1155
rect -5775 1075 -5770 1155
rect -5800 1065 -5770 1075
rect -5710 1155 -5680 1165
rect -5710 1075 -5705 1155
rect -5685 1075 -5680 1155
rect -5710 1065 -5680 1075
rect -5620 1155 -5590 1165
rect -5620 1075 -5615 1155
rect -5595 1075 -5590 1155
rect -5620 1065 -5590 1075
rect -5530 1155 -5500 1165
rect -5530 1075 -5525 1155
rect -5505 1075 -5500 1155
rect -5530 1065 -5500 1075
rect -5440 1155 -5410 1165
rect -5440 1075 -5435 1155
rect -5415 1075 -5410 1155
rect -5440 1065 -5410 1075
rect -5350 1155 -5320 1165
rect -5350 1075 -5345 1155
rect -5325 1075 -5320 1155
rect -5350 1065 -5320 1075
rect -5260 1155 -5230 1165
rect -5260 1075 -5255 1155
rect -5235 1075 -5230 1155
rect -5260 1065 -5230 1075
rect -5170 1155 -5140 1165
rect -5170 1075 -5165 1155
rect -5145 1075 -5140 1155
rect -5170 1065 -5140 1075
rect -5080 1155 -5050 1165
rect -5080 1075 -5075 1155
rect -5055 1075 -5050 1155
rect -5080 1065 -5050 1075
rect -4990 1155 -4960 1165
rect -4990 1075 -4985 1155
rect -4965 1075 -4960 1155
rect -4990 1065 -4960 1075
rect -4900 1155 -4870 1165
rect -4900 1075 -4895 1155
rect -4875 1075 -4870 1155
rect -4900 1065 -4870 1075
rect -4810 1155 -4780 1165
rect -4810 1075 -4805 1155
rect -4785 1075 -4780 1155
rect -4810 1065 -4780 1075
rect -4720 1155 -4690 1165
rect -4720 1075 -4715 1155
rect -4695 1075 -4690 1155
rect -4720 1065 -4690 1075
rect -4630 1155 -4600 1165
rect -4630 1075 -4625 1155
rect -4605 1075 -4600 1155
rect -4630 1065 -4600 1075
rect -4540 1155 -4510 1165
rect -4540 1075 -4535 1155
rect -4515 1075 -4510 1155
rect -4540 1065 -4510 1075
rect -4450 1155 -4420 1165
rect -4450 1075 -4445 1155
rect -4425 1075 -4420 1155
rect -4450 1065 -4420 1075
rect -4360 1155 -4330 1165
rect -4360 1075 -4355 1155
rect -4335 1075 -4330 1155
rect -4360 1065 -4330 1075
rect -4270 1155 -4240 1165
rect -4270 1075 -4265 1155
rect -4245 1075 -4240 1155
rect -4270 1065 -4240 1075
rect -4180 1155 -4150 1165
rect -4180 1075 -4175 1155
rect -4155 1075 -4150 1155
rect -4180 1065 -4150 1075
rect -4090 1155 -4060 1165
rect -4090 1075 -4085 1155
rect -4065 1075 -4060 1155
rect -4090 1065 -4060 1075
rect -4000 1155 -3970 1165
rect -4000 1075 -3995 1155
rect -3975 1075 -3970 1155
rect -4000 1065 -3970 1075
rect -3910 1155 -3880 1165
rect -3910 1075 -3905 1155
rect -3885 1075 -3880 1155
rect -3910 1065 -3880 1075
rect -3820 1155 -3790 1165
rect -3820 1075 -3815 1155
rect -3795 1075 -3790 1155
rect -3820 1065 -3790 1075
rect -3730 1155 -3700 1165
rect -3730 1075 -3725 1155
rect -3705 1075 -3700 1155
rect -3730 1065 -3700 1075
rect -3640 1155 -3610 1165
rect -3640 1075 -3635 1155
rect -3615 1075 -3610 1155
rect -3640 1065 -3610 1075
rect -3550 1155 -3520 1165
rect -3550 1075 -3545 1155
rect -3525 1075 -3520 1155
rect -3550 1065 -3520 1075
rect -3460 1155 -3430 1165
rect -3460 1075 -3455 1155
rect -3435 1075 -3430 1155
rect -3460 1065 -3430 1075
rect -3370 1155 -3340 1165
rect -3370 1075 -3365 1155
rect -3345 1075 -3340 1155
rect -3370 1065 -3340 1075
rect -3280 1155 -3250 1165
rect -3280 1075 -3275 1155
rect -3255 1075 -3250 1155
rect -3280 1065 -3250 1075
rect -3190 1155 -3160 1165
rect -3190 1075 -3185 1155
rect -3165 1075 -3160 1155
rect -3190 1065 -3160 1075
rect -3100 1155 -3070 1165
rect -3100 1075 -3095 1155
rect -3075 1075 -3070 1155
rect -3100 1065 -3070 1075
rect -3010 1155 -2980 1165
rect -3010 1075 -3005 1155
rect -2985 1075 -2980 1155
rect -3010 1065 -2980 1075
rect -2920 1155 -2890 1165
rect -2920 1075 -2915 1155
rect -2895 1075 -2890 1155
rect -2920 1065 -2890 1075
rect -2830 1155 -2800 1165
rect -2830 1075 -2825 1155
rect -2805 1075 -2800 1155
rect -2830 1065 -2800 1075
rect -2740 1155 -2710 1165
rect -2740 1075 -2735 1155
rect -2715 1075 -2710 1155
rect -2740 1065 -2710 1075
rect -2650 1155 -2620 1165
rect -2650 1075 -2645 1155
rect -2625 1075 -2620 1155
rect -2650 1065 -2620 1075
rect -2560 1155 -2530 1165
rect -2560 1075 -2555 1155
rect -2535 1075 -2530 1155
rect -2560 1065 -2530 1075
rect -2470 1155 -2440 1165
rect -2470 1075 -2465 1155
rect -2445 1075 -2440 1155
rect -2470 1065 -2440 1075
rect -2380 1155 -2350 1165
rect -2380 1075 -2375 1155
rect -2355 1075 -2350 1155
rect -2380 1065 -2350 1075
rect -2290 1155 -2260 1165
rect -2290 1075 -2285 1155
rect -2265 1075 -2260 1155
rect -2290 1065 -2260 1075
rect -2200 1155 -2170 1165
rect -2200 1075 -2195 1155
rect -2175 1075 -2170 1155
rect -2200 1065 -2170 1075
rect -2110 1155 -2080 1165
rect -2110 1075 -2105 1155
rect -2085 1075 -2080 1155
rect -2110 1065 -2080 1075
rect -2020 1155 -1990 1165
rect -2020 1075 -2015 1155
rect -1995 1075 -1990 1155
rect -2020 1065 -1990 1075
rect -1930 1155 -1900 1165
rect -1930 1075 -1925 1155
rect -1905 1075 -1900 1155
rect -1930 1065 -1900 1075
rect -1840 1155 -1810 1165
rect -1840 1075 -1835 1155
rect -1815 1075 -1810 1155
rect -1840 1065 -1810 1075
rect -1750 1155 -1720 1165
rect -1750 1075 -1745 1155
rect -1725 1075 -1720 1155
rect -1750 1065 -1720 1075
rect -1660 1155 -1630 1165
rect -1660 1075 -1655 1155
rect -1635 1075 -1630 1155
rect -1660 1065 -1630 1075
rect -1570 1155 -1540 1165
rect -1570 1075 -1565 1155
rect -1545 1075 -1540 1155
rect -1570 1065 -1540 1075
rect -1480 1155 -1450 1165
rect -1480 1075 -1475 1155
rect -1455 1075 -1450 1155
rect -1480 1065 -1450 1075
rect -1390 1155 -1360 1165
rect -1390 1075 -1385 1155
rect -1365 1075 -1360 1155
rect -1390 1065 -1360 1075
rect -1300 1155 -1270 1165
rect -1300 1075 -1295 1155
rect -1275 1075 -1270 1155
rect -1300 1065 -1270 1075
rect -1210 1155 -1180 1165
rect -1210 1075 -1205 1155
rect -1185 1075 -1180 1155
rect -1210 1065 -1180 1075
rect -1120 1155 -1090 1165
rect -1120 1075 -1115 1155
rect -1095 1075 -1090 1155
rect -1120 1065 -1090 1075
rect -1030 1155 -1000 1165
rect -1030 1075 -1025 1155
rect -1005 1075 -1000 1155
rect -1030 1065 -1000 1075
rect -940 1155 -910 1165
rect -940 1075 -935 1155
rect -915 1075 -910 1155
rect -940 1065 -910 1075
rect -850 1155 -820 1165
rect -850 1075 -845 1155
rect -825 1075 -820 1155
rect -850 1065 -820 1075
rect -760 1155 -730 1165
rect -760 1075 -755 1155
rect -735 1075 -730 1155
rect -760 1065 -730 1075
rect -670 1065 -640 1165
rect -580 1065 -550 1165
rect -490 1065 -460 1165
rect -400 1065 -370 1165
rect -310 1065 -280 1165
rect -220 1065 -190 1165
rect -130 1065 -100 1165
rect -40 1155 -10 1165
rect -40 1075 -35 1155
rect -15 1075 -10 1155
rect -40 1065 -10 1075
rect -11555 1045 -11535 1065
rect -11565 1040 -11525 1045
rect -11565 1010 -11560 1040
rect -11530 1010 -11525 1040
rect -11565 1005 -11525 1010
rect -11565 985 -11525 990
rect -11565 955 -11560 985
rect -11530 955 -11525 985
rect -11565 950 -11525 955
rect -11555 930 -11535 950
rect -11465 930 -11445 1065
rect -11375 930 -11355 1065
rect -11285 930 -11265 1065
rect -11195 930 -11175 1065
rect -11105 930 -11085 1065
rect -11015 930 -10995 1065
rect -10925 930 -10905 1065
rect -10835 1045 -10815 1065
rect -9395 1045 -9375 1065
rect -7955 1045 -7935 1065
rect -4355 1045 -4335 1065
rect -755 1045 -735 1065
rect -10845 1040 -10805 1045
rect -10845 1010 -10840 1040
rect -10810 1010 -10805 1040
rect -10845 1005 -10805 1010
rect -10665 1040 -10625 1045
rect -10665 1010 -10660 1040
rect -10630 1010 -10625 1040
rect -10665 1005 -10625 1010
rect -10485 1040 -10445 1045
rect -10485 1010 -10480 1040
rect -10450 1010 -10445 1040
rect -10485 1005 -10445 1010
rect -10305 1040 -10265 1045
rect -10305 1010 -10300 1040
rect -10270 1010 -10265 1040
rect -10305 1005 -10265 1010
rect -10125 1040 -10085 1045
rect -10125 1010 -10120 1040
rect -10090 1010 -10085 1040
rect -10125 1005 -10085 1010
rect -9945 1040 -9905 1045
rect -9945 1010 -9940 1040
rect -9910 1010 -9905 1040
rect -9945 1005 -9905 1010
rect -9765 1040 -9725 1045
rect -9765 1010 -9760 1040
rect -9730 1010 -9725 1040
rect -9765 1005 -9725 1010
rect -9585 1040 -9545 1045
rect -9585 1010 -9580 1040
rect -9550 1010 -9545 1040
rect -9585 1005 -9545 1010
rect -9405 1040 -9365 1045
rect -9405 1010 -9400 1040
rect -9370 1010 -9365 1040
rect -9405 1005 -9365 1010
rect -9225 1040 -9185 1045
rect -9225 1010 -9220 1040
rect -9190 1010 -9185 1040
rect -9225 1005 -9185 1010
rect -9045 1040 -9005 1045
rect -9045 1010 -9040 1040
rect -9010 1010 -9005 1040
rect -9045 1005 -9005 1010
rect -8865 1040 -8825 1045
rect -8865 1010 -8860 1040
rect -8830 1010 -8825 1040
rect -8865 1005 -8825 1010
rect -8685 1040 -8645 1045
rect -8685 1010 -8680 1040
rect -8650 1010 -8645 1040
rect -8685 1005 -8645 1010
rect -8505 1040 -8465 1045
rect -8505 1010 -8500 1040
rect -8470 1010 -8465 1040
rect -8505 1005 -8465 1010
rect -8325 1040 -8285 1045
rect -8325 1010 -8320 1040
rect -8290 1010 -8285 1040
rect -8325 1005 -8285 1010
rect -8145 1040 -8105 1045
rect -8145 1010 -8140 1040
rect -8110 1010 -8105 1040
rect -8145 1005 -8105 1010
rect -7965 1040 -7925 1045
rect -7965 1010 -7960 1040
rect -7930 1010 -7925 1040
rect -7965 1005 -7925 1010
rect -7785 1040 -7745 1045
rect -7785 1010 -7780 1040
rect -7750 1010 -7745 1040
rect -7785 1005 -7745 1010
rect -7605 1040 -7565 1045
rect -7605 1010 -7600 1040
rect -7570 1010 -7565 1040
rect -7605 1005 -7565 1010
rect -7425 1040 -7385 1045
rect -7425 1010 -7420 1040
rect -7390 1010 -7385 1040
rect -7425 1005 -7385 1010
rect -7245 1040 -7205 1045
rect -7245 1010 -7240 1040
rect -7210 1010 -7205 1040
rect -7245 1005 -7205 1010
rect -7065 1040 -7025 1045
rect -7065 1010 -7060 1040
rect -7030 1010 -7025 1040
rect -7065 1005 -7025 1010
rect -6885 1040 -6845 1045
rect -6885 1010 -6880 1040
rect -6850 1010 -6845 1040
rect -6885 1005 -6845 1010
rect -6705 1040 -6665 1045
rect -6705 1010 -6700 1040
rect -6670 1010 -6665 1040
rect -6705 1005 -6665 1010
rect -6525 1040 -6485 1045
rect -6525 1010 -6520 1040
rect -6490 1010 -6485 1040
rect -6525 1005 -6485 1010
rect -6345 1040 -6305 1045
rect -6345 1010 -6340 1040
rect -6310 1010 -6305 1040
rect -6345 1005 -6305 1010
rect -6165 1040 -6125 1045
rect -6165 1010 -6160 1040
rect -6130 1010 -6125 1040
rect -6165 1005 -6125 1010
rect -5985 1040 -5945 1045
rect -5985 1010 -5980 1040
rect -5950 1010 -5945 1040
rect -5985 1005 -5945 1010
rect -5805 1040 -5765 1045
rect -5805 1010 -5800 1040
rect -5770 1010 -5765 1040
rect -5805 1005 -5765 1010
rect -5625 1040 -5585 1045
rect -5625 1010 -5620 1040
rect -5590 1010 -5585 1040
rect -5625 1005 -5585 1010
rect -5445 1040 -5405 1045
rect -5445 1010 -5440 1040
rect -5410 1010 -5405 1040
rect -5445 1005 -5405 1010
rect -5265 1040 -5225 1045
rect -5265 1010 -5260 1040
rect -5230 1010 -5225 1040
rect -5265 1005 -5225 1010
rect -5085 1040 -5045 1045
rect -5085 1010 -5080 1040
rect -5050 1010 -5045 1040
rect -5085 1005 -5045 1010
rect -4905 1040 -4865 1045
rect -4905 1010 -4900 1040
rect -4870 1010 -4865 1040
rect -4905 1005 -4865 1010
rect -4725 1040 -4685 1045
rect -4725 1010 -4720 1040
rect -4690 1010 -4685 1040
rect -4725 1005 -4685 1010
rect -4545 1040 -4505 1045
rect -4545 1010 -4540 1040
rect -4510 1010 -4505 1040
rect -4545 1005 -4505 1010
rect -4365 1040 -4325 1045
rect -4365 1010 -4360 1040
rect -4330 1010 -4325 1040
rect -4365 1005 -4325 1010
rect -4185 1040 -4145 1045
rect -4185 1010 -4180 1040
rect -4150 1010 -4145 1040
rect -4185 1005 -4145 1010
rect -4005 1040 -3965 1045
rect -4005 1010 -4000 1040
rect -3970 1010 -3965 1040
rect -4005 1005 -3965 1010
rect -3825 1040 -3785 1045
rect -3825 1010 -3820 1040
rect -3790 1010 -3785 1040
rect -3825 1005 -3785 1010
rect -3645 1040 -3605 1045
rect -3645 1010 -3640 1040
rect -3610 1010 -3605 1040
rect -3645 1005 -3605 1010
rect -3465 1040 -3425 1045
rect -3465 1010 -3460 1040
rect -3430 1010 -3425 1040
rect -3465 1005 -3425 1010
rect -3285 1040 -3245 1045
rect -3285 1010 -3280 1040
rect -3250 1010 -3245 1040
rect -3285 1005 -3245 1010
rect -3105 1040 -3065 1045
rect -3105 1010 -3100 1040
rect -3070 1010 -3065 1040
rect -3105 1005 -3065 1010
rect -2925 1040 -2885 1045
rect -2925 1010 -2920 1040
rect -2890 1010 -2885 1040
rect -2925 1005 -2885 1010
rect -2745 1040 -2705 1045
rect -2745 1010 -2740 1040
rect -2710 1010 -2705 1040
rect -2745 1005 -2705 1010
rect -2565 1040 -2525 1045
rect -2565 1010 -2560 1040
rect -2530 1010 -2525 1040
rect -2565 1005 -2525 1010
rect -2385 1040 -2345 1045
rect -2385 1010 -2380 1040
rect -2350 1010 -2345 1040
rect -2385 1005 -2345 1010
rect -2205 1040 -2165 1045
rect -2205 1010 -2200 1040
rect -2170 1010 -2165 1040
rect -2205 1005 -2165 1010
rect -2025 1040 -1985 1045
rect -2025 1010 -2020 1040
rect -1990 1010 -1985 1040
rect -2025 1005 -1985 1010
rect -1845 1040 -1805 1045
rect -1845 1010 -1840 1040
rect -1810 1010 -1805 1040
rect -1845 1005 -1805 1010
rect -1665 1040 -1625 1045
rect -1665 1010 -1660 1040
rect -1630 1010 -1625 1040
rect -1665 1005 -1625 1010
rect -1485 1040 -1445 1045
rect -1485 1010 -1480 1040
rect -1450 1010 -1445 1040
rect -1485 1005 -1445 1010
rect -1305 1040 -1265 1045
rect -1305 1010 -1300 1040
rect -1270 1010 -1265 1040
rect -1305 1005 -1265 1010
rect -1125 1040 -1085 1045
rect -1125 1010 -1120 1040
rect -1090 1010 -1085 1040
rect -1125 1005 -1085 1010
rect -945 1040 -905 1045
rect -945 1010 -940 1040
rect -910 1010 -905 1040
rect -945 1005 -905 1010
rect -765 1040 -725 1045
rect -765 1010 -760 1040
rect -730 1010 -725 1040
rect -765 1005 -725 1010
rect -10845 985 -10805 990
rect -10845 955 -10840 985
rect -10810 955 -10805 985
rect -10845 950 -10805 955
rect -10665 985 -10625 990
rect -10665 955 -10660 985
rect -10630 955 -10625 985
rect -10665 950 -10625 955
rect -10485 985 -10445 990
rect -10485 955 -10480 985
rect -10450 955 -10445 985
rect -10485 950 -10445 955
rect -10305 985 -10265 990
rect -10305 955 -10300 985
rect -10270 955 -10265 985
rect -10305 950 -10265 955
rect -10125 985 -10085 990
rect -10125 955 -10120 985
rect -10090 955 -10085 985
rect -10125 950 -10085 955
rect -9945 985 -9905 990
rect -9945 955 -9940 985
rect -9910 955 -9905 985
rect -9945 950 -9905 955
rect -9765 985 -9725 990
rect -9765 955 -9760 985
rect -9730 955 -9725 985
rect -9765 950 -9725 955
rect -9585 985 -9545 990
rect -9585 955 -9580 985
rect -9550 955 -9545 985
rect -9585 950 -9545 955
rect -9405 985 -9365 990
rect -9405 955 -9400 985
rect -9370 955 -9365 985
rect -9405 950 -9365 955
rect -9225 985 -9185 990
rect -9225 955 -9220 985
rect -9190 955 -9185 985
rect -9225 950 -9185 955
rect -9045 985 -9005 990
rect -9045 955 -9040 985
rect -9010 955 -9005 985
rect -9045 950 -9005 955
rect -8865 985 -8825 990
rect -8865 955 -8860 985
rect -8830 955 -8825 985
rect -8865 950 -8825 955
rect -8685 985 -8645 990
rect -8685 955 -8680 985
rect -8650 955 -8645 985
rect -8685 950 -8645 955
rect -8505 985 -8465 990
rect -8505 955 -8500 985
rect -8470 955 -8465 985
rect -8505 950 -8465 955
rect -8325 985 -8285 990
rect -8325 955 -8320 985
rect -8290 955 -8285 985
rect -8325 950 -8285 955
rect -8145 985 -8105 990
rect -8145 955 -8140 985
rect -8110 955 -8105 985
rect -8145 950 -8105 955
rect -7965 985 -7925 990
rect -7965 955 -7960 985
rect -7930 955 -7925 985
rect -7965 950 -7925 955
rect -7785 985 -7745 990
rect -7785 955 -7780 985
rect -7750 955 -7745 985
rect -7785 950 -7745 955
rect -7605 985 -7565 990
rect -7605 955 -7600 985
rect -7570 955 -7565 985
rect -7605 950 -7565 955
rect -7425 985 -7385 990
rect -7425 955 -7420 985
rect -7390 955 -7385 985
rect -7425 950 -7385 955
rect -7245 985 -7205 990
rect -7245 955 -7240 985
rect -7210 955 -7205 985
rect -7245 950 -7205 955
rect -7065 985 -7025 990
rect -7065 955 -7060 985
rect -7030 955 -7025 985
rect -7065 950 -7025 955
rect -6885 985 -6845 990
rect -6885 955 -6880 985
rect -6850 955 -6845 985
rect -6885 950 -6845 955
rect -6705 985 -6665 990
rect -6705 955 -6700 985
rect -6670 955 -6665 985
rect -6705 950 -6665 955
rect -6525 985 -6485 990
rect -6525 955 -6520 985
rect -6490 955 -6485 985
rect -6525 950 -6485 955
rect -6345 985 -6305 990
rect -6345 955 -6340 985
rect -6310 955 -6305 985
rect -6345 950 -6305 955
rect -6165 985 -6125 990
rect -6165 955 -6160 985
rect -6130 955 -6125 985
rect -6165 950 -6125 955
rect -5985 985 -5945 990
rect -5985 955 -5980 985
rect -5950 955 -5945 985
rect -5985 950 -5945 955
rect -5805 985 -5765 990
rect -5805 955 -5800 985
rect -5770 955 -5765 985
rect -5805 950 -5765 955
rect -5625 985 -5585 990
rect -5625 955 -5620 985
rect -5590 955 -5585 985
rect -5625 950 -5585 955
rect -5445 985 -5405 990
rect -5445 955 -5440 985
rect -5410 955 -5405 985
rect -5445 950 -5405 955
rect -5265 985 -5225 990
rect -5265 955 -5260 985
rect -5230 955 -5225 985
rect -5265 950 -5225 955
rect -5085 985 -5045 990
rect -5085 955 -5080 985
rect -5050 955 -5045 985
rect -5085 950 -5045 955
rect -4905 985 -4865 990
rect -4905 955 -4900 985
rect -4870 955 -4865 985
rect -4905 950 -4865 955
rect -4725 985 -4685 990
rect -4725 955 -4720 985
rect -4690 955 -4685 985
rect -4725 950 -4685 955
rect -4545 985 -4505 990
rect -4545 955 -4540 985
rect -4510 955 -4505 985
rect -4545 950 -4505 955
rect -4365 985 -4325 990
rect -4365 955 -4360 985
rect -4330 955 -4325 985
rect -4365 950 -4325 955
rect -4185 985 -4145 990
rect -4185 955 -4180 985
rect -4150 955 -4145 985
rect -4185 950 -4145 955
rect -4005 985 -3965 990
rect -4005 955 -4000 985
rect -3970 955 -3965 985
rect -4005 950 -3965 955
rect -3825 985 -3785 990
rect -3825 955 -3820 985
rect -3790 955 -3785 985
rect -3825 950 -3785 955
rect -3645 985 -3605 990
rect -3645 955 -3640 985
rect -3610 955 -3605 985
rect -3645 950 -3605 955
rect -3465 985 -3425 990
rect -3465 955 -3460 985
rect -3430 955 -3425 985
rect -3465 950 -3425 955
rect -3285 985 -3245 990
rect -3285 955 -3280 985
rect -3250 955 -3245 985
rect -3285 950 -3245 955
rect -3105 985 -3065 990
rect -3105 955 -3100 985
rect -3070 955 -3065 985
rect -3105 950 -3065 955
rect -2925 985 -2885 990
rect -2925 955 -2920 985
rect -2890 955 -2885 985
rect -2925 950 -2885 955
rect -2745 985 -2705 990
rect -2745 955 -2740 985
rect -2710 955 -2705 985
rect -2745 950 -2705 955
rect -2565 985 -2525 990
rect -2565 955 -2560 985
rect -2530 955 -2525 985
rect -2565 950 -2525 955
rect -2385 985 -2345 990
rect -2385 955 -2380 985
rect -2350 955 -2345 985
rect -2385 950 -2345 955
rect -2205 985 -2165 990
rect -2205 955 -2200 985
rect -2170 955 -2165 985
rect -2205 950 -2165 955
rect -2025 985 -1985 990
rect -2025 955 -2020 985
rect -1990 955 -1985 985
rect -2025 950 -1985 955
rect -1845 985 -1805 990
rect -1845 955 -1840 985
rect -1810 955 -1805 985
rect -1845 950 -1805 955
rect -1665 985 -1625 990
rect -1665 955 -1660 985
rect -1630 955 -1625 985
rect -1665 950 -1625 955
rect -1485 985 -1445 990
rect -1485 955 -1480 985
rect -1450 955 -1445 985
rect -1485 950 -1445 955
rect -1305 985 -1265 990
rect -1305 955 -1300 985
rect -1270 955 -1265 985
rect -1305 950 -1265 955
rect -1125 985 -1085 990
rect -1125 955 -1120 985
rect -1090 955 -1085 985
rect -1125 950 -1085 955
rect -945 985 -905 990
rect -945 955 -940 985
rect -910 955 -905 985
rect -945 950 -905 955
rect -765 985 -725 990
rect -765 955 -760 985
rect -730 955 -725 985
rect -765 950 -725 955
rect -10835 930 -10815 950
rect -7235 930 -7215 950
rect -3635 930 -3615 950
rect -2195 930 -2175 950
rect -755 930 -735 950
rect -665 930 -645 1065
rect -575 930 -555 1065
rect -485 930 -465 1065
rect -395 930 -375 1065
rect -305 930 -285 1065
rect -215 930 -195 1065
rect -125 930 -105 1065
rect -35 1045 -15 1065
rect -45 1040 -5 1045
rect -45 1010 -40 1040
rect -10 1010 -5 1040
rect -45 1005 -5 1010
rect -45 985 -5 990
rect -45 955 -40 985
rect -10 955 -5 985
rect -45 950 -5 955
rect -35 930 -15 950
rect -11560 920 -11530 930
rect -11560 840 -11555 920
rect -11535 840 -11530 920
rect -11560 830 -11530 840
rect -11470 830 -11440 930
rect -11380 830 -11350 930
rect -11290 830 -11260 930
rect -11200 830 -11170 930
rect -11110 830 -11080 930
rect -11020 830 -10990 930
rect -10930 830 -10900 930
rect -10840 920 -10810 930
rect -10840 840 -10835 920
rect -10815 840 -10810 920
rect -10840 830 -10810 840
rect -10750 920 -10720 930
rect -10750 840 -10745 920
rect -10725 840 -10720 920
rect -10750 830 -10720 840
rect -10660 920 -10630 930
rect -10660 840 -10655 920
rect -10635 840 -10630 920
rect -10660 830 -10630 840
rect -10570 920 -10540 930
rect -10570 840 -10565 920
rect -10545 840 -10540 920
rect -10570 830 -10540 840
rect -10480 920 -10450 930
rect -10480 840 -10475 920
rect -10455 840 -10450 920
rect -10480 830 -10450 840
rect -10390 920 -10360 930
rect -10390 840 -10385 920
rect -10365 840 -10360 920
rect -10390 830 -10360 840
rect -10300 920 -10270 930
rect -10300 840 -10295 920
rect -10275 840 -10270 920
rect -10300 830 -10270 840
rect -10210 920 -10180 930
rect -10210 840 -10205 920
rect -10185 840 -10180 920
rect -10210 830 -10180 840
rect -10120 920 -10090 930
rect -10120 840 -10115 920
rect -10095 840 -10090 920
rect -10120 830 -10090 840
rect -10030 920 -10000 930
rect -10030 840 -10025 920
rect -10005 840 -10000 920
rect -10030 830 -10000 840
rect -9940 920 -9910 930
rect -9940 840 -9935 920
rect -9915 840 -9910 920
rect -9940 830 -9910 840
rect -9850 920 -9820 930
rect -9850 840 -9845 920
rect -9825 840 -9820 920
rect -9850 830 -9820 840
rect -9760 920 -9730 930
rect -9760 840 -9755 920
rect -9735 840 -9730 920
rect -9760 830 -9730 840
rect -9670 920 -9640 930
rect -9670 840 -9665 920
rect -9645 840 -9640 920
rect -9670 830 -9640 840
rect -9580 920 -9550 930
rect -9580 840 -9575 920
rect -9555 840 -9550 920
rect -9580 830 -9550 840
rect -9490 920 -9460 930
rect -9490 840 -9485 920
rect -9465 840 -9460 920
rect -9490 830 -9460 840
rect -9400 920 -9370 930
rect -9400 840 -9395 920
rect -9375 840 -9370 920
rect -9400 830 -9370 840
rect -9310 920 -9280 930
rect -9310 840 -9305 920
rect -9285 840 -9280 920
rect -9310 830 -9280 840
rect -9220 920 -9190 930
rect -9220 840 -9215 920
rect -9195 840 -9190 920
rect -9220 830 -9190 840
rect -9130 920 -9100 930
rect -9130 840 -9125 920
rect -9105 840 -9100 920
rect -9130 830 -9100 840
rect -9040 920 -9010 930
rect -9040 840 -9035 920
rect -9015 840 -9010 920
rect -9040 830 -9010 840
rect -8950 920 -8920 930
rect -8950 840 -8945 920
rect -8925 840 -8920 920
rect -8950 830 -8920 840
rect -8860 920 -8830 930
rect -8860 840 -8855 920
rect -8835 840 -8830 920
rect -8860 830 -8830 840
rect -8770 920 -8740 930
rect -8770 840 -8765 920
rect -8745 840 -8740 920
rect -8770 830 -8740 840
rect -8680 920 -8650 930
rect -8680 840 -8675 920
rect -8655 840 -8650 920
rect -8680 830 -8650 840
rect -8590 920 -8560 930
rect -8590 840 -8585 920
rect -8565 840 -8560 920
rect -8590 830 -8560 840
rect -8500 920 -8470 930
rect -8500 840 -8495 920
rect -8475 840 -8470 920
rect -8500 830 -8470 840
rect -8410 920 -8380 930
rect -8410 840 -8405 920
rect -8385 840 -8380 920
rect -8410 830 -8380 840
rect -8320 920 -8290 930
rect -8320 840 -8315 920
rect -8295 840 -8290 920
rect -8320 830 -8290 840
rect -8230 920 -8200 930
rect -8230 840 -8225 920
rect -8205 840 -8200 920
rect -8230 830 -8200 840
rect -8140 920 -8110 930
rect -8140 840 -8135 920
rect -8115 840 -8110 920
rect -8140 830 -8110 840
rect -8050 920 -8020 930
rect -8050 840 -8045 920
rect -8025 840 -8020 920
rect -8050 830 -8020 840
rect -7960 920 -7930 930
rect -7960 840 -7955 920
rect -7935 840 -7930 920
rect -7960 830 -7930 840
rect -7870 920 -7840 930
rect -7870 840 -7865 920
rect -7845 840 -7840 920
rect -7870 830 -7840 840
rect -7780 920 -7750 930
rect -7780 840 -7775 920
rect -7755 840 -7750 920
rect -7780 830 -7750 840
rect -7690 920 -7660 930
rect -7690 840 -7685 920
rect -7665 840 -7660 920
rect -7690 830 -7660 840
rect -7600 920 -7570 930
rect -7600 840 -7595 920
rect -7575 840 -7570 920
rect -7600 830 -7570 840
rect -7510 920 -7480 930
rect -7510 840 -7505 920
rect -7485 840 -7480 920
rect -7510 830 -7480 840
rect -7420 920 -7390 930
rect -7420 840 -7415 920
rect -7395 840 -7390 920
rect -7420 830 -7390 840
rect -7330 920 -7300 930
rect -7330 840 -7325 920
rect -7305 840 -7300 920
rect -7330 830 -7300 840
rect -7240 920 -7210 930
rect -7240 840 -7235 920
rect -7215 840 -7210 920
rect -7240 830 -7210 840
rect -7150 920 -7120 930
rect -7150 840 -7145 920
rect -7125 840 -7120 920
rect -7150 830 -7120 840
rect -7060 920 -7030 930
rect -7060 840 -7055 920
rect -7035 840 -7030 920
rect -7060 830 -7030 840
rect -6970 920 -6940 930
rect -6970 840 -6965 920
rect -6945 840 -6940 920
rect -6970 830 -6940 840
rect -6880 920 -6850 930
rect -6880 840 -6875 920
rect -6855 840 -6850 920
rect -6880 830 -6850 840
rect -6790 920 -6760 930
rect -6790 840 -6785 920
rect -6765 840 -6760 920
rect -6790 830 -6760 840
rect -6700 920 -6670 930
rect -6700 840 -6695 920
rect -6675 840 -6670 920
rect -6700 830 -6670 840
rect -6610 920 -6580 930
rect -6610 840 -6605 920
rect -6585 840 -6580 920
rect -6610 830 -6580 840
rect -6520 920 -6490 930
rect -6520 840 -6515 920
rect -6495 840 -6490 920
rect -6520 830 -6490 840
rect -6430 920 -6400 930
rect -6430 840 -6425 920
rect -6405 840 -6400 920
rect -6430 830 -6400 840
rect -6340 920 -6310 930
rect -6340 840 -6335 920
rect -6315 840 -6310 920
rect -6340 830 -6310 840
rect -6250 920 -6220 930
rect -6250 840 -6245 920
rect -6225 840 -6220 920
rect -6250 830 -6220 840
rect -6160 920 -6130 930
rect -6160 840 -6155 920
rect -6135 840 -6130 920
rect -6160 830 -6130 840
rect -6070 920 -6040 930
rect -6070 840 -6065 920
rect -6045 840 -6040 920
rect -6070 830 -6040 840
rect -5980 920 -5950 930
rect -5980 840 -5975 920
rect -5955 840 -5950 920
rect -5980 830 -5950 840
rect -5890 920 -5860 930
rect -5890 840 -5885 920
rect -5865 840 -5860 920
rect -5890 830 -5860 840
rect -5800 920 -5770 930
rect -5800 840 -5795 920
rect -5775 840 -5770 920
rect -5800 830 -5770 840
rect -5710 920 -5680 930
rect -5710 840 -5705 920
rect -5685 840 -5680 920
rect -5710 830 -5680 840
rect -5620 920 -5590 930
rect -5620 840 -5615 920
rect -5595 840 -5590 920
rect -5620 830 -5590 840
rect -5530 920 -5500 930
rect -5530 840 -5525 920
rect -5505 840 -5500 920
rect -5530 830 -5500 840
rect -5440 920 -5410 930
rect -5440 840 -5435 920
rect -5415 840 -5410 920
rect -5440 830 -5410 840
rect -5350 920 -5320 930
rect -5350 840 -5345 920
rect -5325 840 -5320 920
rect -5350 830 -5320 840
rect -5260 920 -5230 930
rect -5260 840 -5255 920
rect -5235 840 -5230 920
rect -5260 830 -5230 840
rect -5170 920 -5140 930
rect -5170 840 -5165 920
rect -5145 840 -5140 920
rect -5170 830 -5140 840
rect -5080 920 -5050 930
rect -5080 840 -5075 920
rect -5055 840 -5050 920
rect -5080 830 -5050 840
rect -4990 920 -4960 930
rect -4990 840 -4985 920
rect -4965 840 -4960 920
rect -4990 830 -4960 840
rect -4900 920 -4870 930
rect -4900 840 -4895 920
rect -4875 840 -4870 920
rect -4900 830 -4870 840
rect -4810 920 -4780 930
rect -4810 840 -4805 920
rect -4785 840 -4780 920
rect -4810 830 -4780 840
rect -4720 920 -4690 930
rect -4720 840 -4715 920
rect -4695 840 -4690 920
rect -4720 830 -4690 840
rect -4630 920 -4600 930
rect -4630 840 -4625 920
rect -4605 840 -4600 920
rect -4630 830 -4600 840
rect -4540 920 -4510 930
rect -4540 840 -4535 920
rect -4515 840 -4510 920
rect -4540 830 -4510 840
rect -4450 920 -4420 930
rect -4450 840 -4445 920
rect -4425 840 -4420 920
rect -4450 830 -4420 840
rect -4360 920 -4330 930
rect -4360 840 -4355 920
rect -4335 840 -4330 920
rect -4360 830 -4330 840
rect -4270 920 -4240 930
rect -4270 840 -4265 920
rect -4245 840 -4240 920
rect -4270 830 -4240 840
rect -4180 920 -4150 930
rect -4180 840 -4175 920
rect -4155 840 -4150 920
rect -4180 830 -4150 840
rect -4090 920 -4060 930
rect -4090 840 -4085 920
rect -4065 840 -4060 920
rect -4090 830 -4060 840
rect -4000 920 -3970 930
rect -4000 840 -3995 920
rect -3975 840 -3970 920
rect -4000 830 -3970 840
rect -3910 920 -3880 930
rect -3910 840 -3905 920
rect -3885 840 -3880 920
rect -3910 830 -3880 840
rect -3820 920 -3790 930
rect -3820 840 -3815 920
rect -3795 840 -3790 920
rect -3820 830 -3790 840
rect -3730 920 -3700 930
rect -3730 840 -3725 920
rect -3705 840 -3700 920
rect -3730 830 -3700 840
rect -3640 920 -3610 930
rect -3640 840 -3635 920
rect -3615 840 -3610 920
rect -3640 830 -3610 840
rect -3550 920 -3520 930
rect -3550 840 -3545 920
rect -3525 840 -3520 920
rect -3550 830 -3520 840
rect -3460 920 -3430 930
rect -3460 840 -3455 920
rect -3435 840 -3430 920
rect -3460 830 -3430 840
rect -3370 920 -3340 930
rect -3370 840 -3365 920
rect -3345 840 -3340 920
rect -3370 830 -3340 840
rect -3280 920 -3250 930
rect -3280 840 -3275 920
rect -3255 840 -3250 920
rect -3280 830 -3250 840
rect -3190 920 -3160 930
rect -3190 840 -3185 920
rect -3165 840 -3160 920
rect -3190 830 -3160 840
rect -3100 920 -3070 930
rect -3100 840 -3095 920
rect -3075 840 -3070 920
rect -3100 830 -3070 840
rect -3010 920 -2980 930
rect -3010 840 -3005 920
rect -2985 840 -2980 920
rect -3010 830 -2980 840
rect -2920 920 -2890 930
rect -2920 840 -2915 920
rect -2895 840 -2890 920
rect -2920 830 -2890 840
rect -2830 920 -2800 930
rect -2830 840 -2825 920
rect -2805 840 -2800 920
rect -2830 830 -2800 840
rect -2740 920 -2710 930
rect -2740 840 -2735 920
rect -2715 840 -2710 920
rect -2740 830 -2710 840
rect -2650 920 -2620 930
rect -2650 840 -2645 920
rect -2625 840 -2620 920
rect -2650 830 -2620 840
rect -2560 920 -2530 930
rect -2560 840 -2555 920
rect -2535 840 -2530 920
rect -2560 830 -2530 840
rect -2470 920 -2440 930
rect -2470 840 -2465 920
rect -2445 840 -2440 920
rect -2470 830 -2440 840
rect -2380 920 -2350 930
rect -2380 840 -2375 920
rect -2355 840 -2350 920
rect -2380 830 -2350 840
rect -2290 920 -2260 930
rect -2290 840 -2285 920
rect -2265 840 -2260 920
rect -2290 830 -2260 840
rect -2200 920 -2170 930
rect -2200 840 -2195 920
rect -2175 840 -2170 920
rect -2200 830 -2170 840
rect -2110 920 -2080 930
rect -2110 840 -2105 920
rect -2085 840 -2080 920
rect -2110 830 -2080 840
rect -2020 920 -1990 930
rect -2020 840 -2015 920
rect -1995 840 -1990 920
rect -2020 830 -1990 840
rect -1930 920 -1900 930
rect -1930 840 -1925 920
rect -1905 840 -1900 920
rect -1930 830 -1900 840
rect -1840 920 -1810 930
rect -1840 840 -1835 920
rect -1815 840 -1810 920
rect -1840 830 -1810 840
rect -1750 920 -1720 930
rect -1750 840 -1745 920
rect -1725 840 -1720 920
rect -1750 830 -1720 840
rect -1660 920 -1630 930
rect -1660 840 -1655 920
rect -1635 840 -1630 920
rect -1660 830 -1630 840
rect -1570 920 -1540 930
rect -1570 840 -1565 920
rect -1545 840 -1540 920
rect -1570 830 -1540 840
rect -1480 920 -1450 930
rect -1480 840 -1475 920
rect -1455 840 -1450 920
rect -1480 830 -1450 840
rect -1390 920 -1360 930
rect -1390 840 -1385 920
rect -1365 840 -1360 920
rect -1390 830 -1360 840
rect -1300 920 -1270 930
rect -1300 840 -1295 920
rect -1275 840 -1270 920
rect -1300 830 -1270 840
rect -1210 920 -1180 930
rect -1210 840 -1205 920
rect -1185 840 -1180 920
rect -1210 830 -1180 840
rect -1120 920 -1090 930
rect -1120 840 -1115 920
rect -1095 840 -1090 920
rect -1120 830 -1090 840
rect -1030 920 -1000 930
rect -1030 840 -1025 920
rect -1005 840 -1000 920
rect -1030 830 -1000 840
rect -940 920 -910 930
rect -940 840 -935 920
rect -915 840 -910 920
rect -940 830 -910 840
rect -850 920 -820 930
rect -850 840 -845 920
rect -825 840 -820 920
rect -850 830 -820 840
rect -760 920 -730 930
rect -760 840 -755 920
rect -735 840 -730 920
rect -760 830 -730 840
rect -670 830 -640 930
rect -580 830 -550 930
rect -490 830 -460 930
rect -400 830 -370 930
rect -310 830 -280 930
rect -220 830 -190 930
rect -130 830 -100 930
rect -40 920 -10 930
rect -40 840 -35 920
rect -15 840 -10 920
rect -40 830 -10 840
rect -11465 525 -11445 830
rect -11470 520 -11440 525
rect -11470 500 -11465 520
rect -11445 500 -11440 520
rect -11470 495 -11440 500
rect -11465 150 -11445 495
rect -11375 485 -11355 830
rect -11380 480 -11350 485
rect -11380 460 -11375 480
rect -11355 460 -11350 480
rect -11380 455 -11350 460
rect -11375 150 -11355 455
rect -11285 445 -11265 830
rect -11290 440 -11260 445
rect -11290 420 -11285 440
rect -11265 420 -11260 440
rect -11290 415 -11260 420
rect -11285 150 -11265 415
rect -11195 405 -11175 830
rect -11200 400 -11170 405
rect -11200 380 -11195 400
rect -11175 380 -11170 400
rect -11200 375 -11170 380
rect -11195 150 -11175 375
rect -11105 365 -11085 830
rect -11110 360 -11080 365
rect -11110 340 -11105 360
rect -11085 340 -11080 360
rect -11110 335 -11080 340
rect -11105 150 -11085 335
rect -11015 150 -10995 830
rect -10925 150 -10905 830
rect -10700 810 -10680 815
rect -10520 810 -10500 815
rect -10340 810 -10320 815
rect -10160 810 -10140 815
rect -10705 805 -10675 810
rect -10705 785 -10700 805
rect -10680 785 -10675 805
rect -10705 780 -10675 785
rect -10525 805 -10495 810
rect -10525 785 -10520 805
rect -10500 785 -10495 805
rect -10525 780 -10495 785
rect -10345 805 -10315 810
rect -10345 785 -10340 805
rect -10320 785 -10315 805
rect -10345 780 -10315 785
rect -10165 805 -10135 810
rect -10165 785 -10160 805
rect -10140 785 -10135 805
rect -10165 780 -10135 785
rect -10700 645 -10680 780
rect -10520 645 -10500 780
rect -10705 640 -10675 645
rect -10705 620 -10700 640
rect -10680 620 -10675 640
rect -10705 615 -10675 620
rect -10525 640 -10495 645
rect -10525 620 -10520 640
rect -10500 620 -10495 640
rect -10525 615 -10495 620
rect -10700 610 -10680 615
rect -10520 610 -10500 615
rect -10340 605 -10320 780
rect -10160 605 -10140 780
rect -10115 725 -10095 830
rect -10120 720 -10090 725
rect -10120 700 -10115 720
rect -10095 700 -10090 720
rect -10120 695 -10090 700
rect -10115 690 -10095 695
rect -10345 600 -10315 605
rect -10345 580 -10340 600
rect -10320 580 -10315 600
rect -10345 575 -10315 580
rect -10165 600 -10135 605
rect -10165 580 -10160 600
rect -10140 580 -10135 600
rect -10165 575 -10135 580
rect -10340 570 -10320 575
rect -10160 570 -10140 575
rect -10115 565 -10095 570
rect -10120 560 -10090 565
rect -10120 540 -10115 560
rect -10095 540 -10090 560
rect -10120 535 -10090 540
rect -10475 365 -10455 370
rect -10480 360 -10450 365
rect -10480 340 -10475 360
rect -10455 340 -10450 360
rect -10480 335 -10450 340
rect -10790 285 -10770 290
rect -10610 285 -10590 290
rect -10795 280 -10765 285
rect -10795 260 -10790 280
rect -10770 260 -10765 280
rect -10795 255 -10765 260
rect -10615 280 -10585 285
rect -10615 260 -10610 280
rect -10590 260 -10585 280
rect -10615 255 -10585 260
rect -10790 200 -10770 255
rect -10610 200 -10590 255
rect -10795 195 -10765 200
rect -10795 175 -10790 195
rect -10770 175 -10765 195
rect -10795 170 -10765 175
rect -10615 195 -10585 200
rect -10615 175 -10610 195
rect -10590 175 -10585 195
rect -10615 170 -10585 175
rect -10790 165 -10770 170
rect -10610 165 -10590 170
rect -10475 150 -10455 335
rect -10430 325 -10410 330
rect -10250 325 -10230 330
rect -10435 320 -10405 325
rect -10435 300 -10430 320
rect -10410 300 -10405 320
rect -10435 295 -10405 300
rect -10255 320 -10225 325
rect -10255 300 -10250 320
rect -10230 300 -10225 320
rect -10255 295 -10225 300
rect -10430 200 -10410 295
rect -10250 200 -10230 295
rect -10435 195 -10405 200
rect -10435 175 -10430 195
rect -10410 175 -10405 195
rect -10435 170 -10405 175
rect -10255 195 -10225 200
rect -10255 175 -10250 195
rect -10230 175 -10225 195
rect -10255 170 -10225 175
rect -10430 165 -10410 170
rect -10250 165 -10230 170
rect -10115 150 -10095 535
rect -10025 365 -10005 830
rect -9980 810 -9960 815
rect -9985 805 -9955 810
rect -9985 785 -9980 805
rect -9960 785 -9955 805
rect -9985 780 -9955 785
rect -9980 445 -9960 780
rect -9935 725 -9915 830
rect -9940 720 -9910 725
rect -9940 700 -9935 720
rect -9915 700 -9910 720
rect -9940 695 -9910 700
rect -9935 690 -9915 695
rect -9985 440 -9955 445
rect -9985 420 -9980 440
rect -9960 420 -9955 440
rect -9985 415 -9955 420
rect -9980 410 -9960 415
rect -9845 365 -9825 830
rect -9800 810 -9780 815
rect -9805 805 -9775 810
rect -9805 785 -9800 805
rect -9780 785 -9775 805
rect -9805 780 -9775 785
rect -9800 445 -9780 780
rect -9755 725 -9735 830
rect -9760 720 -9730 725
rect -9760 700 -9755 720
rect -9735 700 -9730 720
rect -9760 695 -9730 700
rect -9755 690 -9735 695
rect -9805 440 -9775 445
rect -9805 420 -9800 440
rect -9780 420 -9775 440
rect -9805 415 -9775 420
rect -9800 410 -9780 415
rect -9665 365 -9645 830
rect -9620 810 -9600 815
rect -9625 805 -9595 810
rect -9625 785 -9620 805
rect -9600 785 -9595 805
rect -9625 780 -9595 785
rect -9620 445 -9600 780
rect -9575 725 -9555 830
rect -9580 720 -9550 725
rect -9580 700 -9575 720
rect -9555 700 -9550 720
rect -9580 695 -9550 700
rect -9575 690 -9555 695
rect -9625 440 -9595 445
rect -9625 420 -9620 440
rect -9600 420 -9595 440
rect -9625 415 -9595 420
rect -9620 410 -9600 415
rect -9485 365 -9465 830
rect -9440 810 -9420 815
rect -9445 805 -9415 810
rect -9445 785 -9440 805
rect -9420 785 -9415 805
rect -9445 780 -9415 785
rect -9440 445 -9420 780
rect -9395 725 -9375 830
rect -9400 720 -9370 725
rect -9400 700 -9395 720
rect -9375 700 -9370 720
rect -9400 695 -9370 700
rect -9395 690 -9375 695
rect -9445 440 -9415 445
rect -9445 420 -9440 440
rect -9420 420 -9415 440
rect -9445 415 -9415 420
rect -9440 410 -9420 415
rect -9305 365 -9285 830
rect -9260 810 -9240 815
rect -9265 805 -9235 810
rect -9265 785 -9260 805
rect -9240 785 -9235 805
rect -9265 780 -9235 785
rect -9260 445 -9240 780
rect -9215 725 -9195 830
rect -9220 720 -9190 725
rect -9220 700 -9215 720
rect -9195 700 -9190 720
rect -9220 695 -9190 700
rect -9215 690 -9195 695
rect -9265 440 -9235 445
rect -9265 420 -9260 440
rect -9240 420 -9235 440
rect -9265 415 -9235 420
rect -9260 410 -9240 415
rect -9125 365 -9105 830
rect -9080 810 -9060 815
rect -9085 805 -9055 810
rect -9085 785 -9080 805
rect -9060 785 -9055 805
rect -9085 780 -9055 785
rect -9080 445 -9060 780
rect -9035 725 -9015 830
rect -9040 720 -9010 725
rect -9040 700 -9035 720
rect -9015 700 -9010 720
rect -9040 695 -9010 700
rect -9035 690 -9015 695
rect -9085 440 -9055 445
rect -9085 420 -9080 440
rect -9060 420 -9055 440
rect -9085 415 -9055 420
rect -9080 410 -9060 415
rect -8945 365 -8925 830
rect -8900 810 -8880 815
rect -8905 805 -8875 810
rect -8905 785 -8900 805
rect -8880 785 -8875 805
rect -8905 780 -8875 785
rect -8900 445 -8880 780
rect -8855 725 -8835 830
rect -8860 720 -8830 725
rect -8860 700 -8855 720
rect -8835 700 -8830 720
rect -8860 695 -8830 700
rect -8855 690 -8835 695
rect -8905 440 -8875 445
rect -8905 420 -8900 440
rect -8880 420 -8875 440
rect -8905 415 -8875 420
rect -8900 410 -8880 415
rect -8765 365 -8745 830
rect -8720 810 -8700 815
rect -8725 805 -8695 810
rect -8725 785 -8720 805
rect -8700 785 -8695 805
rect -8725 780 -8695 785
rect -8720 445 -8700 780
rect -8675 725 -8655 830
rect -8680 720 -8650 725
rect -8680 700 -8675 720
rect -8655 700 -8650 720
rect -8680 695 -8650 700
rect -8675 690 -8655 695
rect -8725 440 -8695 445
rect -8725 420 -8720 440
rect -8700 420 -8695 440
rect -8725 415 -8695 420
rect -8720 410 -8700 415
rect -8585 365 -8565 830
rect -8540 810 -8520 815
rect -8545 805 -8515 810
rect -8545 785 -8540 805
rect -8520 785 -8515 805
rect -8545 780 -8515 785
rect -8540 445 -8520 780
rect -8495 725 -8475 830
rect -8500 720 -8470 725
rect -8500 700 -8495 720
rect -8475 700 -8470 720
rect -8500 695 -8470 700
rect -8495 690 -8475 695
rect -8545 440 -8515 445
rect -8545 420 -8540 440
rect -8520 420 -8515 440
rect -8545 415 -8515 420
rect -8540 410 -8520 415
rect -8405 365 -8385 830
rect -8360 810 -8340 815
rect -8365 805 -8335 810
rect -8365 785 -8360 805
rect -8340 785 -8335 805
rect -8365 780 -8335 785
rect -8360 445 -8340 780
rect -8315 725 -8295 830
rect -8320 720 -8290 725
rect -8320 700 -8315 720
rect -8295 700 -8290 720
rect -8320 695 -8290 700
rect -8315 690 -8295 695
rect -8365 440 -8335 445
rect -8365 420 -8360 440
rect -8340 420 -8335 440
rect -8365 415 -8335 420
rect -8360 410 -8340 415
rect -8225 365 -8205 830
rect -8180 810 -8160 815
rect -8185 805 -8155 810
rect -8185 785 -8180 805
rect -8160 785 -8155 805
rect -8185 780 -8155 785
rect -8180 445 -8160 780
rect -8135 725 -8115 830
rect -8140 720 -8110 725
rect -8140 700 -8135 720
rect -8115 700 -8110 720
rect -8140 695 -8110 700
rect -8135 690 -8115 695
rect -8185 440 -8155 445
rect -8185 420 -8180 440
rect -8160 420 -8155 440
rect -8185 415 -8155 420
rect -8180 410 -8160 415
rect -8045 365 -8025 830
rect -8000 810 -7980 815
rect -8005 805 -7975 810
rect -8005 785 -8000 805
rect -7980 785 -7975 805
rect -8005 780 -7975 785
rect -8000 445 -7980 780
rect -7955 725 -7935 830
rect -7820 810 -7800 815
rect -7640 810 -7620 815
rect -7460 810 -7440 815
rect -7280 810 -7260 815
rect -7100 810 -7080 815
rect -6920 810 -6900 815
rect -6740 810 -6720 815
rect -6560 810 -6540 815
rect -7825 805 -7795 810
rect -7825 785 -7820 805
rect -7800 785 -7795 805
rect -7825 780 -7795 785
rect -7645 805 -7615 810
rect -7645 785 -7640 805
rect -7620 785 -7615 805
rect -7645 780 -7615 785
rect -7465 805 -7435 810
rect -7465 785 -7460 805
rect -7440 785 -7435 805
rect -7465 780 -7435 785
rect -7285 805 -7255 810
rect -7285 785 -7280 805
rect -7260 785 -7255 805
rect -7285 780 -7255 785
rect -7105 805 -7075 810
rect -7105 785 -7100 805
rect -7080 785 -7075 805
rect -7105 780 -7075 785
rect -6925 805 -6895 810
rect -6925 785 -6920 805
rect -6900 785 -6895 805
rect -6925 780 -6895 785
rect -6745 805 -6715 810
rect -6745 785 -6740 805
rect -6720 785 -6715 805
rect -6745 780 -6715 785
rect -6565 805 -6535 810
rect -6565 785 -6560 805
rect -6540 785 -6535 805
rect -6565 780 -6535 785
rect -7960 720 -7930 725
rect -7960 700 -7955 720
rect -7935 700 -7930 720
rect -7960 695 -7930 700
rect -7955 690 -7935 695
rect -7820 605 -7800 780
rect -7640 605 -7620 780
rect -7460 645 -7440 780
rect -7280 645 -7260 780
rect -7100 645 -7080 780
rect -6920 645 -6900 780
rect -7465 640 -7435 645
rect -7465 620 -7460 640
rect -7440 620 -7435 640
rect -7465 615 -7435 620
rect -7285 640 -7255 645
rect -7285 620 -7280 640
rect -7260 620 -7255 640
rect -7285 615 -7255 620
rect -7105 640 -7075 645
rect -7105 620 -7100 640
rect -7080 620 -7075 640
rect -7105 615 -7075 620
rect -6925 640 -6895 645
rect -6925 620 -6920 640
rect -6900 620 -6895 640
rect -6925 615 -6895 620
rect -7460 610 -7440 615
rect -7280 610 -7260 615
rect -7100 610 -7080 615
rect -6920 610 -6900 615
rect -6740 605 -6720 780
rect -6560 605 -6540 780
rect -6515 725 -6495 830
rect -6520 720 -6490 725
rect -6520 700 -6515 720
rect -6495 700 -6490 720
rect -6520 695 -6490 700
rect -6515 690 -6495 695
rect -7825 600 -7795 605
rect -7825 580 -7820 600
rect -7800 580 -7795 600
rect -7825 575 -7795 580
rect -7645 600 -7615 605
rect -7645 580 -7640 600
rect -7620 580 -7615 600
rect -7645 575 -7615 580
rect -6745 600 -6715 605
rect -6745 580 -6740 600
rect -6720 580 -6715 600
rect -6745 575 -6715 580
rect -6565 600 -6535 605
rect -6565 580 -6560 600
rect -6540 580 -6535 600
rect -6565 575 -6535 580
rect -7820 570 -7800 575
rect -7640 570 -7620 575
rect -6740 570 -6720 575
rect -6560 570 -6540 575
rect -7955 565 -7935 570
rect -7960 560 -7930 565
rect -7960 540 -7955 560
rect -7935 540 -7930 560
rect -7960 535 -7930 540
rect -8005 440 -7975 445
rect -8005 420 -8000 440
rect -7980 420 -7975 440
rect -8005 415 -7975 420
rect -8000 410 -7980 415
rect -10030 360 -10000 365
rect -10030 340 -10025 360
rect -10005 340 -10000 360
rect -10030 335 -10000 340
rect -9850 360 -9820 365
rect -9850 340 -9845 360
rect -9825 340 -9820 360
rect -9850 335 -9820 340
rect -9670 360 -9640 365
rect -9670 340 -9665 360
rect -9645 340 -9640 360
rect -9670 335 -9640 340
rect -9490 360 -9460 365
rect -9490 340 -9485 360
rect -9465 340 -9460 360
rect -9490 335 -9460 340
rect -9310 360 -9280 365
rect -9310 340 -9305 360
rect -9285 340 -9280 360
rect -9310 335 -9280 340
rect -9130 360 -9100 365
rect -9130 340 -9125 360
rect -9105 340 -9100 360
rect -9130 335 -9100 340
rect -8950 360 -8920 365
rect -8950 340 -8945 360
rect -8925 340 -8920 360
rect -8950 335 -8920 340
rect -8770 360 -8740 365
rect -8770 340 -8765 360
rect -8745 340 -8740 360
rect -8770 335 -8740 340
rect -8590 360 -8560 365
rect -8590 340 -8585 360
rect -8565 340 -8560 360
rect -8590 335 -8560 340
rect -8410 360 -8380 365
rect -8410 340 -8405 360
rect -8385 340 -8380 360
rect -8410 335 -8380 340
rect -8230 360 -8200 365
rect -8230 340 -8225 360
rect -8205 340 -8200 360
rect -8230 335 -8200 340
rect -8050 360 -8020 365
rect -8050 340 -8045 360
rect -8025 340 -8020 360
rect -8050 335 -8020 340
rect -10025 330 -10005 335
rect -9845 330 -9825 335
rect -9665 330 -9645 335
rect -9485 330 -9465 335
rect -9305 330 -9285 335
rect -9125 330 -9105 335
rect -8945 330 -8925 335
rect -8765 330 -8745 335
rect -8585 330 -8565 335
rect -8405 330 -8385 335
rect -8225 330 -8205 335
rect -8045 330 -8025 335
rect -10070 200 -10050 205
rect -9890 200 -9870 205
rect -9710 200 -9690 205
rect -9530 200 -9510 205
rect -9350 200 -9330 205
rect -9170 200 -9150 205
rect -8990 200 -8970 205
rect -8810 200 -8790 205
rect -8630 200 -8610 205
rect -8450 200 -8430 205
rect -8270 200 -8250 205
rect -8090 200 -8070 205
rect -10075 195 -10045 200
rect -10075 175 -10070 195
rect -10050 175 -10045 195
rect -10075 170 -10045 175
rect -9895 195 -9865 200
rect -9895 175 -9890 195
rect -9870 175 -9865 195
rect -9895 170 -9865 175
rect -9715 195 -9685 200
rect -9715 175 -9710 195
rect -9690 175 -9685 195
rect -9715 170 -9685 175
rect -9535 195 -9505 200
rect -9535 175 -9530 195
rect -9510 175 -9505 195
rect -9535 170 -9505 175
rect -9355 195 -9325 200
rect -9355 175 -9350 195
rect -9330 175 -9325 195
rect -9355 170 -9325 175
rect -9175 195 -9145 200
rect -9175 175 -9170 195
rect -9150 175 -9145 195
rect -9175 170 -9145 175
rect -8995 195 -8965 200
rect -8995 175 -8990 195
rect -8970 175 -8965 195
rect -8995 170 -8965 175
rect -8815 195 -8785 200
rect -8815 175 -8810 195
rect -8790 175 -8785 195
rect -8815 170 -8785 175
rect -8635 195 -8605 200
rect -8635 175 -8630 195
rect -8610 175 -8605 195
rect -8635 170 -8605 175
rect -8455 195 -8425 200
rect -8455 175 -8450 195
rect -8430 175 -8425 195
rect -8455 170 -8425 175
rect -8275 195 -8245 200
rect -8275 175 -8270 195
rect -8250 175 -8245 195
rect -8275 170 -8245 175
rect -8095 195 -8065 200
rect -8095 175 -8090 195
rect -8070 175 -8065 195
rect -8095 170 -8065 175
rect -10070 165 -10050 170
rect -9890 165 -9870 170
rect -9710 165 -9690 170
rect -9530 165 -9510 170
rect -9350 165 -9330 170
rect -9170 165 -9150 170
rect -8990 165 -8970 170
rect -8810 165 -8790 170
rect -8630 165 -8610 170
rect -8450 165 -8430 170
rect -8270 165 -8250 170
rect -8090 165 -8070 170
rect -7955 150 -7935 535
rect -6515 525 -6495 530
rect -6520 520 -6490 525
rect -6520 500 -6515 520
rect -6495 500 -6490 520
rect -6520 495 -6490 500
rect -6875 405 -6855 410
rect -6880 400 -6850 405
rect -6880 380 -6875 400
rect -6855 380 -6850 400
rect -6880 375 -6850 380
rect -7595 365 -7575 370
rect -7600 360 -7570 365
rect -7600 340 -7595 360
rect -7575 340 -7570 360
rect -7600 335 -7570 340
rect -7910 325 -7890 330
rect -7730 325 -7710 330
rect -7915 320 -7885 325
rect -7915 300 -7910 320
rect -7890 300 -7885 320
rect -7915 295 -7885 300
rect -7735 320 -7705 325
rect -7735 300 -7730 320
rect -7710 300 -7705 320
rect -7735 295 -7705 300
rect -7910 200 -7890 295
rect -7730 200 -7710 295
rect -7915 195 -7885 200
rect -7915 175 -7910 195
rect -7890 175 -7885 195
rect -7915 170 -7885 175
rect -7735 195 -7705 200
rect -7735 175 -7730 195
rect -7710 175 -7705 195
rect -7735 170 -7705 175
rect -7910 165 -7890 170
rect -7730 165 -7710 170
rect -7595 150 -7575 335
rect -7550 285 -7530 290
rect -7370 285 -7350 290
rect -7190 285 -7170 290
rect -7010 285 -6990 290
rect -7555 280 -7525 285
rect -7555 260 -7550 280
rect -7530 260 -7525 280
rect -7555 255 -7525 260
rect -7375 280 -7345 285
rect -7375 260 -7370 280
rect -7350 260 -7345 280
rect -7375 255 -7345 260
rect -7195 280 -7165 285
rect -7195 260 -7190 280
rect -7170 260 -7165 280
rect -7195 255 -7165 260
rect -7015 280 -6985 285
rect -7015 260 -7010 280
rect -6990 260 -6985 280
rect -7015 255 -6985 260
rect -7550 200 -7530 255
rect -7370 200 -7350 255
rect -7190 200 -7170 255
rect -7010 200 -6990 255
rect -7555 195 -7525 200
rect -7555 175 -7550 195
rect -7530 175 -7525 195
rect -7555 170 -7525 175
rect -7375 195 -7345 200
rect -7375 175 -7370 195
rect -7350 175 -7345 195
rect -7375 170 -7345 175
rect -7195 195 -7165 200
rect -7195 175 -7190 195
rect -7170 175 -7165 195
rect -7195 170 -7165 175
rect -7015 195 -6985 200
rect -7015 175 -7010 195
rect -6990 175 -6985 195
rect -7015 170 -6985 175
rect -7550 165 -7530 170
rect -7370 165 -7350 170
rect -7190 165 -7170 170
rect -7010 165 -6990 170
rect -6875 150 -6855 375
rect -6830 325 -6810 330
rect -6650 325 -6630 330
rect -6835 320 -6805 325
rect -6835 300 -6830 320
rect -6810 300 -6805 320
rect -6835 295 -6805 300
rect -6655 320 -6625 325
rect -6655 300 -6650 320
rect -6630 300 -6625 320
rect -6655 295 -6625 300
rect -6830 200 -6810 295
rect -6650 200 -6630 295
rect -6835 195 -6805 200
rect -6835 175 -6830 195
rect -6810 175 -6805 195
rect -6835 170 -6805 175
rect -6655 195 -6625 200
rect -6655 175 -6650 195
rect -6630 175 -6625 195
rect -6655 170 -6625 175
rect -6830 165 -6810 170
rect -6650 165 -6630 170
rect -6515 150 -6495 495
rect -6425 405 -6405 830
rect -6380 810 -6360 815
rect -6385 805 -6355 810
rect -6385 785 -6380 805
rect -6360 785 -6355 805
rect -6385 780 -6355 785
rect -6380 485 -6360 780
rect -6335 725 -6315 830
rect -6340 720 -6310 725
rect -6340 700 -6335 720
rect -6315 700 -6310 720
rect -6340 695 -6310 700
rect -6335 690 -6315 695
rect -6385 480 -6355 485
rect -6385 460 -6380 480
rect -6360 460 -6355 480
rect -6385 455 -6355 460
rect -6380 450 -6360 455
rect -6245 405 -6225 830
rect -6200 810 -6180 815
rect -6205 805 -6175 810
rect -6205 785 -6200 805
rect -6180 785 -6175 805
rect -6205 780 -6175 785
rect -6200 485 -6180 780
rect -6155 725 -6135 830
rect -6160 720 -6130 725
rect -6160 700 -6155 720
rect -6135 700 -6130 720
rect -6160 695 -6130 700
rect -6155 690 -6135 695
rect -6205 480 -6175 485
rect -6205 460 -6200 480
rect -6180 460 -6175 480
rect -6205 455 -6175 460
rect -6200 450 -6180 455
rect -6065 405 -6045 830
rect -6020 810 -6000 815
rect -6025 805 -5995 810
rect -6025 785 -6020 805
rect -6000 785 -5995 805
rect -6025 780 -5995 785
rect -6020 485 -6000 780
rect -5975 725 -5955 830
rect -5980 720 -5950 725
rect -5980 700 -5975 720
rect -5955 700 -5950 720
rect -5980 695 -5950 700
rect -5975 690 -5955 695
rect -6025 480 -5995 485
rect -6025 460 -6020 480
rect -6000 460 -5995 480
rect -6025 455 -5995 460
rect -6020 450 -6000 455
rect -5885 405 -5865 830
rect -5840 810 -5820 815
rect -5845 805 -5815 810
rect -5845 785 -5840 805
rect -5820 785 -5815 805
rect -5845 780 -5815 785
rect -5840 485 -5820 780
rect -5795 725 -5775 830
rect -5800 720 -5770 725
rect -5800 700 -5795 720
rect -5775 700 -5770 720
rect -5800 695 -5770 700
rect -5795 690 -5775 695
rect -5845 480 -5815 485
rect -5845 460 -5840 480
rect -5820 460 -5815 480
rect -5845 455 -5815 460
rect -5840 450 -5820 455
rect -5705 405 -5685 830
rect -5660 810 -5640 815
rect -5665 805 -5635 810
rect -5665 785 -5660 805
rect -5640 785 -5635 805
rect -5665 780 -5635 785
rect -5660 485 -5640 780
rect -5615 725 -5595 830
rect -5620 720 -5590 725
rect -5620 700 -5615 720
rect -5595 700 -5590 720
rect -5620 695 -5590 700
rect -5615 690 -5595 695
rect -5665 480 -5635 485
rect -5665 460 -5660 480
rect -5640 460 -5635 480
rect -5665 455 -5635 460
rect -5660 450 -5640 455
rect -5525 405 -5505 830
rect -5480 810 -5460 815
rect -5485 805 -5455 810
rect -5485 785 -5480 805
rect -5460 785 -5455 805
rect -5485 780 -5455 785
rect -5480 485 -5460 780
rect -5435 725 -5415 830
rect -5440 720 -5410 725
rect -5440 700 -5435 720
rect -5415 700 -5410 720
rect -5440 695 -5410 700
rect -5435 690 -5415 695
rect -5485 480 -5455 485
rect -5485 460 -5480 480
rect -5460 460 -5455 480
rect -5485 455 -5455 460
rect -5480 450 -5460 455
rect -5345 405 -5325 830
rect -5300 810 -5280 815
rect -5305 805 -5275 810
rect -5305 785 -5300 805
rect -5280 785 -5275 805
rect -5305 780 -5275 785
rect -5300 485 -5280 780
rect -5255 725 -5235 830
rect -5260 720 -5230 725
rect -5260 700 -5255 720
rect -5235 700 -5230 720
rect -5260 695 -5230 700
rect -5255 690 -5235 695
rect -5305 480 -5275 485
rect -5305 460 -5300 480
rect -5280 460 -5275 480
rect -5305 455 -5275 460
rect -5300 450 -5280 455
rect -5165 405 -5145 830
rect -5120 810 -5100 815
rect -5125 805 -5095 810
rect -5125 785 -5120 805
rect -5100 785 -5095 805
rect -5125 780 -5095 785
rect -5120 485 -5100 780
rect -5075 725 -5055 830
rect -5080 720 -5050 725
rect -5080 700 -5075 720
rect -5055 700 -5050 720
rect -5080 695 -5050 700
rect -5075 690 -5055 695
rect -5125 480 -5095 485
rect -5125 460 -5120 480
rect -5100 460 -5095 480
rect -5125 455 -5095 460
rect -5120 450 -5100 455
rect -4985 405 -4965 830
rect -4940 810 -4920 815
rect -4945 805 -4915 810
rect -4945 785 -4940 805
rect -4920 785 -4915 805
rect -4945 780 -4915 785
rect -4940 485 -4920 780
rect -4895 725 -4875 830
rect -4900 720 -4870 725
rect -4900 700 -4895 720
rect -4875 700 -4870 720
rect -4900 695 -4870 700
rect -4895 690 -4875 695
rect -4945 480 -4915 485
rect -4945 460 -4940 480
rect -4920 460 -4915 480
rect -4945 455 -4915 460
rect -4940 450 -4920 455
rect -4805 405 -4785 830
rect -4760 810 -4740 815
rect -4765 805 -4735 810
rect -4765 785 -4760 805
rect -4740 785 -4735 805
rect -4765 780 -4735 785
rect -4760 485 -4740 780
rect -4715 725 -4695 830
rect -4720 720 -4690 725
rect -4720 700 -4715 720
rect -4695 700 -4690 720
rect -4720 695 -4690 700
rect -4715 690 -4695 695
rect -4765 480 -4735 485
rect -4765 460 -4760 480
rect -4740 460 -4735 480
rect -4765 455 -4735 460
rect -4760 450 -4740 455
rect -4625 405 -4605 830
rect -4580 810 -4560 815
rect -4585 805 -4555 810
rect -4585 785 -4580 805
rect -4560 785 -4555 805
rect -4585 780 -4555 785
rect -4580 485 -4560 780
rect -4535 725 -4515 830
rect -4540 720 -4510 725
rect -4540 700 -4535 720
rect -4515 700 -4510 720
rect -4540 695 -4510 700
rect -4535 690 -4515 695
rect -4585 480 -4555 485
rect -4585 460 -4580 480
rect -4560 460 -4555 480
rect -4585 455 -4555 460
rect -4580 450 -4560 455
rect -4445 405 -4425 830
rect -4400 810 -4380 815
rect -4405 805 -4375 810
rect -4405 785 -4400 805
rect -4380 785 -4375 805
rect -4405 780 -4375 785
rect -4400 485 -4380 780
rect -4355 725 -4335 830
rect -4220 810 -4200 815
rect -4040 810 -4020 815
rect -3860 810 -3840 815
rect -3680 810 -3660 815
rect -3500 810 -3480 815
rect -3320 810 -3300 815
rect -3140 810 -3120 815
rect -2960 810 -2940 815
rect -4225 805 -4195 810
rect -4225 785 -4220 805
rect -4200 785 -4195 805
rect -4225 780 -4195 785
rect -4045 805 -4015 810
rect -4045 785 -4040 805
rect -4020 785 -4015 805
rect -4045 780 -4015 785
rect -3865 805 -3835 810
rect -3865 785 -3860 805
rect -3840 785 -3835 805
rect -3865 780 -3835 785
rect -3685 805 -3655 810
rect -3685 785 -3680 805
rect -3660 785 -3655 805
rect -3685 780 -3655 785
rect -3505 805 -3475 810
rect -3505 785 -3500 805
rect -3480 785 -3475 805
rect -3505 780 -3475 785
rect -3325 805 -3295 810
rect -3325 785 -3320 805
rect -3300 785 -3295 805
rect -3325 780 -3295 785
rect -3145 805 -3115 810
rect -3145 785 -3140 805
rect -3120 785 -3115 805
rect -3145 780 -3115 785
rect -2965 805 -2935 810
rect -2965 785 -2960 805
rect -2940 785 -2935 805
rect -2965 780 -2935 785
rect -4360 720 -4330 725
rect -4360 700 -4355 720
rect -4335 700 -4330 720
rect -4360 695 -4330 700
rect -4355 690 -4335 695
rect -4220 605 -4200 780
rect -4040 605 -4020 780
rect -3860 645 -3840 780
rect -3680 645 -3660 780
rect -3865 640 -3835 645
rect -3865 620 -3860 640
rect -3840 620 -3835 640
rect -3865 615 -3835 620
rect -3685 640 -3655 645
rect -3685 620 -3680 640
rect -3660 620 -3655 640
rect -3685 615 -3655 620
rect -3860 610 -3840 615
rect -3680 610 -3660 615
rect -4225 600 -4195 605
rect -4225 580 -4220 600
rect -4200 580 -4195 600
rect -4225 575 -4195 580
rect -4045 600 -4015 605
rect -4045 580 -4040 600
rect -4020 580 -4015 600
rect -4045 575 -4015 580
rect -4220 570 -4200 575
rect -4040 570 -4020 575
rect -3500 565 -3480 780
rect -3320 565 -3300 780
rect -3140 605 -3120 780
rect -2960 605 -2940 780
rect -3145 600 -3115 605
rect -3145 580 -3140 600
rect -3120 580 -3115 600
rect -3145 575 -3115 580
rect -2965 600 -2935 605
rect -2965 580 -2960 600
rect -2940 580 -2935 600
rect -2965 575 -2935 580
rect -3140 570 -3120 575
rect -2960 570 -2940 575
rect -2915 565 -2895 830
rect -2780 810 -2760 815
rect -2600 810 -2580 815
rect -2420 810 -2400 815
rect -2240 810 -2220 815
rect -2060 810 -2040 815
rect -1880 810 -1860 815
rect -1700 810 -1680 815
rect -1520 810 -1500 815
rect -2785 805 -2755 810
rect -2785 785 -2780 805
rect -2760 785 -2755 805
rect -2785 780 -2755 785
rect -2605 805 -2575 810
rect -2605 785 -2600 805
rect -2580 785 -2575 805
rect -2605 780 -2575 785
rect -2425 805 -2395 810
rect -2425 785 -2420 805
rect -2400 785 -2395 805
rect -2425 780 -2395 785
rect -2245 805 -2215 810
rect -2245 785 -2240 805
rect -2220 785 -2215 805
rect -2245 780 -2215 785
rect -2065 805 -2035 810
rect -2065 785 -2060 805
rect -2040 785 -2035 805
rect -2065 780 -2035 785
rect -1885 805 -1855 810
rect -1885 785 -1880 805
rect -1860 785 -1855 805
rect -1885 780 -1855 785
rect -1705 805 -1675 810
rect -1705 785 -1700 805
rect -1680 785 -1675 805
rect -1705 780 -1675 785
rect -1525 805 -1495 810
rect -1525 785 -1520 805
rect -1500 785 -1495 805
rect -1525 780 -1495 785
rect -2780 605 -2760 780
rect -2600 605 -2580 780
rect -2785 600 -2755 605
rect -2785 580 -2780 600
rect -2760 580 -2755 600
rect -2785 575 -2755 580
rect -2605 600 -2575 605
rect -2605 580 -2600 600
rect -2580 580 -2575 600
rect -2605 575 -2575 580
rect -2780 570 -2760 575
rect -2600 570 -2580 575
rect -2420 565 -2400 780
rect -2240 565 -2220 780
rect -2060 565 -2040 780
rect -1880 565 -1860 780
rect -1700 605 -1680 780
rect -1520 605 -1500 780
rect -1705 600 -1675 605
rect -1705 580 -1700 600
rect -1680 580 -1675 600
rect -1705 575 -1675 580
rect -1525 600 -1495 605
rect -1525 580 -1520 600
rect -1500 580 -1495 600
rect -1525 575 -1495 580
rect -1700 570 -1680 575
rect -1520 570 -1500 575
rect -3505 560 -3475 565
rect -3505 540 -3500 560
rect -3480 540 -3475 560
rect -3505 535 -3475 540
rect -3325 560 -3295 565
rect -3325 540 -3320 560
rect -3300 540 -3295 560
rect -3325 535 -3295 540
rect -2920 560 -2890 565
rect -2920 540 -2915 560
rect -2895 540 -2890 560
rect -2920 535 -2890 540
rect -2425 560 -2395 565
rect -2425 540 -2420 560
rect -2400 540 -2395 560
rect -2425 535 -2395 540
rect -2245 560 -2215 565
rect -2245 540 -2240 560
rect -2220 540 -2215 560
rect -2245 535 -2215 540
rect -2065 560 -2035 565
rect -2065 540 -2060 560
rect -2040 540 -2035 560
rect -2065 535 -2035 540
rect -1885 560 -1855 565
rect -1885 540 -1880 560
rect -1860 540 -1855 560
rect -1885 535 -1855 540
rect -3500 530 -3480 535
rect -3320 530 -3300 535
rect -4355 525 -4335 530
rect -4360 520 -4330 525
rect -4360 500 -4355 520
rect -4335 500 -4330 520
rect -4360 495 -4330 500
rect -4405 480 -4375 485
rect -4405 460 -4400 480
rect -4380 460 -4375 480
rect -4405 455 -4375 460
rect -4400 450 -4380 455
rect -6430 400 -6400 405
rect -6430 380 -6425 400
rect -6405 380 -6400 400
rect -6430 375 -6400 380
rect -6250 400 -6220 405
rect -6250 380 -6245 400
rect -6225 380 -6220 400
rect -6250 375 -6220 380
rect -6070 400 -6040 405
rect -6070 380 -6065 400
rect -6045 380 -6040 400
rect -6070 375 -6040 380
rect -5890 400 -5860 405
rect -5890 380 -5885 400
rect -5865 380 -5860 400
rect -5890 375 -5860 380
rect -5710 400 -5680 405
rect -5710 380 -5705 400
rect -5685 380 -5680 400
rect -5710 375 -5680 380
rect -5530 400 -5500 405
rect -5530 380 -5525 400
rect -5505 380 -5500 400
rect -5530 375 -5500 380
rect -5350 400 -5320 405
rect -5350 380 -5345 400
rect -5325 380 -5320 400
rect -5350 375 -5320 380
rect -5170 400 -5140 405
rect -5170 380 -5165 400
rect -5145 380 -5140 400
rect -5170 375 -5140 380
rect -4990 400 -4960 405
rect -4990 380 -4985 400
rect -4965 380 -4960 400
rect -4990 375 -4960 380
rect -4810 400 -4780 405
rect -4810 380 -4805 400
rect -4785 380 -4780 400
rect -4810 375 -4780 380
rect -4630 400 -4600 405
rect -4630 380 -4625 400
rect -4605 380 -4600 400
rect -4630 375 -4600 380
rect -4450 400 -4420 405
rect -4450 380 -4445 400
rect -4425 380 -4420 400
rect -4450 375 -4420 380
rect -6425 370 -6405 375
rect -6245 370 -6225 375
rect -6065 370 -6045 375
rect -5885 370 -5865 375
rect -5705 370 -5685 375
rect -5525 370 -5505 375
rect -5345 370 -5325 375
rect -5165 370 -5145 375
rect -4985 370 -4965 375
rect -4805 370 -4785 375
rect -4625 370 -4605 375
rect -4445 370 -4425 375
rect -6470 200 -6450 205
rect -6290 200 -6270 205
rect -6110 200 -6090 205
rect -5930 200 -5910 205
rect -5750 200 -5730 205
rect -5570 200 -5550 205
rect -5390 200 -5370 205
rect -5210 200 -5190 205
rect -5030 200 -5010 205
rect -4850 200 -4830 205
rect -4670 200 -4650 205
rect -4490 200 -4470 205
rect -6475 195 -6445 200
rect -6475 175 -6470 195
rect -6450 175 -6445 195
rect -6475 170 -6445 175
rect -6295 195 -6265 200
rect -6295 175 -6290 195
rect -6270 175 -6265 195
rect -6295 170 -6265 175
rect -6115 195 -6085 200
rect -6115 175 -6110 195
rect -6090 175 -6085 195
rect -6115 170 -6085 175
rect -5935 195 -5905 200
rect -5935 175 -5930 195
rect -5910 175 -5905 195
rect -5935 170 -5905 175
rect -5755 195 -5725 200
rect -5755 175 -5750 195
rect -5730 175 -5725 195
rect -5755 170 -5725 175
rect -5575 195 -5545 200
rect -5575 175 -5570 195
rect -5550 175 -5545 195
rect -5575 170 -5545 175
rect -5395 195 -5365 200
rect -5395 175 -5390 195
rect -5370 175 -5365 195
rect -5395 170 -5365 175
rect -5215 195 -5185 200
rect -5215 175 -5210 195
rect -5190 175 -5185 195
rect -5215 170 -5185 175
rect -5035 195 -5005 200
rect -5035 175 -5030 195
rect -5010 175 -5005 195
rect -5035 170 -5005 175
rect -4855 195 -4825 200
rect -4855 175 -4850 195
rect -4830 175 -4825 195
rect -4855 170 -4825 175
rect -4675 195 -4645 200
rect -4675 175 -4670 195
rect -4650 175 -4645 195
rect -4675 170 -4645 175
rect -4495 195 -4465 200
rect -4495 175 -4490 195
rect -4470 175 -4465 195
rect -4495 170 -4465 175
rect -6470 165 -6450 170
rect -6290 165 -6270 170
rect -6110 165 -6090 170
rect -5930 165 -5910 170
rect -5750 165 -5730 170
rect -5570 165 -5550 170
rect -5390 165 -5370 170
rect -5210 165 -5190 170
rect -5030 165 -5010 170
rect -4850 165 -4830 170
rect -4670 165 -4650 170
rect -4490 165 -4470 170
rect -4355 150 -4335 495
rect -3995 405 -3975 410
rect -4000 400 -3970 405
rect -4000 380 -3995 400
rect -3975 380 -3970 400
rect -4000 375 -3970 380
rect -4310 325 -4290 330
rect -4130 325 -4110 330
rect -4315 320 -4285 325
rect -4315 300 -4310 320
rect -4290 300 -4285 320
rect -4315 295 -4285 300
rect -4135 320 -4105 325
rect -4135 300 -4130 320
rect -4110 300 -4105 320
rect -4135 295 -4105 300
rect -4310 200 -4290 295
rect -4130 200 -4110 295
rect -4315 195 -4285 200
rect -4315 175 -4310 195
rect -4290 175 -4285 195
rect -4315 170 -4285 175
rect -4135 195 -4105 200
rect -4135 175 -4130 195
rect -4110 175 -4105 195
rect -4135 170 -4105 175
rect -4310 165 -4290 170
rect -4130 165 -4110 170
rect -3995 150 -3975 375
rect -3275 365 -3255 370
rect -3280 360 -3250 365
rect -3280 340 -3275 360
rect -3255 340 -3250 360
rect -3280 335 -3250 340
rect -3950 285 -3930 290
rect -3770 285 -3750 290
rect -3590 285 -3570 290
rect -3410 285 -3390 290
rect -3955 280 -3925 285
rect -3955 260 -3950 280
rect -3930 260 -3925 280
rect -3955 255 -3925 260
rect -3775 280 -3745 285
rect -3775 260 -3770 280
rect -3750 260 -3745 280
rect -3775 255 -3745 260
rect -3595 280 -3565 285
rect -3595 260 -3590 280
rect -3570 260 -3565 280
rect -3595 255 -3565 260
rect -3415 280 -3385 285
rect -3415 260 -3410 280
rect -3390 260 -3385 280
rect -3415 255 -3385 260
rect -3950 200 -3930 255
rect -3770 200 -3750 255
rect -3590 200 -3570 255
rect -3410 200 -3390 255
rect -3955 195 -3925 200
rect -3955 175 -3950 195
rect -3930 175 -3925 195
rect -3955 170 -3925 175
rect -3775 195 -3745 200
rect -3775 175 -3770 195
rect -3750 175 -3745 195
rect -3775 170 -3745 175
rect -3595 195 -3565 200
rect -3595 175 -3590 195
rect -3570 175 -3565 195
rect -3595 170 -3565 175
rect -3415 195 -3385 200
rect -3415 175 -3410 195
rect -3390 175 -3385 195
rect -3415 170 -3385 175
rect -3950 165 -3930 170
rect -3770 165 -3750 170
rect -3590 165 -3570 170
rect -3410 165 -3390 170
rect -3275 150 -3255 335
rect -3230 325 -3210 330
rect -3050 325 -3030 330
rect -3235 320 -3205 325
rect -3235 300 -3230 320
rect -3210 300 -3205 320
rect -3235 295 -3205 300
rect -3055 320 -3025 325
rect -3055 300 -3050 320
rect -3030 300 -3025 320
rect -3055 295 -3025 300
rect -3230 200 -3210 295
rect -3050 200 -3030 295
rect -3235 195 -3205 200
rect -3235 175 -3230 195
rect -3210 175 -3205 195
rect -3235 170 -3205 175
rect -3055 195 -3025 200
rect -3055 175 -3050 195
rect -3030 175 -3025 195
rect -3055 170 -3025 175
rect -3230 165 -3210 170
rect -3050 165 -3030 170
rect -2915 150 -2895 535
rect -2420 530 -2400 535
rect -2240 530 -2220 535
rect -2060 530 -2040 535
rect -1880 530 -1860 535
rect -1475 525 -1455 830
rect -1340 810 -1320 815
rect -1160 810 -1140 815
rect -980 810 -960 815
rect -800 810 -780 815
rect -1345 805 -1315 810
rect -1345 785 -1340 805
rect -1320 785 -1315 805
rect -1345 780 -1315 785
rect -1165 805 -1135 810
rect -1165 785 -1160 805
rect -1140 785 -1135 805
rect -1165 780 -1135 785
rect -985 805 -955 810
rect -985 785 -980 805
rect -960 785 -955 805
rect -985 780 -955 785
rect -805 805 -775 810
rect -805 785 -800 805
rect -780 785 -775 805
rect -805 780 -775 785
rect -1340 605 -1320 780
rect -1160 605 -1140 780
rect -1345 600 -1315 605
rect -1345 580 -1340 600
rect -1320 580 -1315 600
rect -1345 575 -1315 580
rect -1165 600 -1135 605
rect -1165 580 -1160 600
rect -1140 580 -1135 600
rect -1165 575 -1135 580
rect -1340 570 -1320 575
rect -1160 570 -1140 575
rect -980 565 -960 780
rect -800 565 -780 780
rect -985 560 -955 565
rect -985 540 -980 560
rect -960 540 -955 560
rect -985 535 -955 540
rect -805 560 -775 565
rect -805 540 -800 560
rect -780 540 -775 560
rect -805 535 -775 540
rect -980 530 -960 535
rect -800 530 -780 535
rect -1480 520 -1450 525
rect -1480 500 -1475 520
rect -1455 500 -1450 520
rect -1480 495 -1450 500
rect -1835 405 -1815 410
rect -1840 400 -1810 405
rect -1840 380 -1835 400
rect -1815 380 -1810 400
rect -1840 375 -1810 380
rect -2555 365 -2535 370
rect -2560 360 -2530 365
rect -2560 340 -2555 360
rect -2535 340 -2530 360
rect -2560 335 -2530 340
rect -2870 325 -2850 330
rect -2690 325 -2670 330
rect -2875 320 -2845 325
rect -2875 300 -2870 320
rect -2850 300 -2845 320
rect -2875 295 -2845 300
rect -2695 320 -2665 325
rect -2695 300 -2690 320
rect -2670 300 -2665 320
rect -2695 295 -2665 300
rect -2870 200 -2850 295
rect -2690 200 -2670 295
rect -2875 195 -2845 200
rect -2875 175 -2870 195
rect -2850 175 -2845 195
rect -2875 170 -2845 175
rect -2695 195 -2665 200
rect -2695 175 -2690 195
rect -2670 175 -2665 195
rect -2695 170 -2665 175
rect -2870 165 -2850 170
rect -2690 165 -2670 170
rect -2555 150 -2535 335
rect -2510 285 -2490 290
rect -2330 285 -2310 290
rect -2150 285 -2130 290
rect -1970 285 -1950 290
rect -2515 280 -2485 285
rect -2515 260 -2510 280
rect -2490 260 -2485 280
rect -2515 255 -2485 260
rect -2335 280 -2305 285
rect -2335 260 -2330 280
rect -2310 260 -2305 280
rect -2335 255 -2305 260
rect -2155 280 -2125 285
rect -2155 260 -2150 280
rect -2130 260 -2125 280
rect -2155 255 -2125 260
rect -1975 280 -1945 285
rect -1975 260 -1970 280
rect -1950 260 -1945 280
rect -1975 255 -1945 260
rect -2510 200 -2490 255
rect -2330 200 -2310 255
rect -2150 200 -2130 255
rect -1970 200 -1950 255
rect -2515 195 -2485 200
rect -2515 175 -2510 195
rect -2490 175 -2485 195
rect -2515 170 -2485 175
rect -2335 195 -2305 200
rect -2335 175 -2330 195
rect -2310 175 -2305 195
rect -2335 170 -2305 175
rect -2155 195 -2125 200
rect -2155 175 -2150 195
rect -2130 175 -2125 195
rect -2155 170 -2125 175
rect -1975 195 -1945 200
rect -1975 175 -1970 195
rect -1950 175 -1945 195
rect -1975 170 -1945 175
rect -2510 165 -2490 170
rect -2330 165 -2310 170
rect -2150 165 -2130 170
rect -1970 165 -1950 170
rect -1835 150 -1815 375
rect -1790 325 -1770 330
rect -1610 325 -1590 330
rect -1795 320 -1765 325
rect -1795 300 -1790 320
rect -1770 300 -1765 320
rect -1795 295 -1765 300
rect -1615 320 -1585 325
rect -1615 300 -1610 320
rect -1590 300 -1585 320
rect -1615 295 -1585 300
rect -1790 200 -1770 295
rect -1610 200 -1590 295
rect -1795 195 -1765 200
rect -1795 175 -1790 195
rect -1770 175 -1765 195
rect -1795 170 -1765 175
rect -1615 195 -1585 200
rect -1615 175 -1610 195
rect -1590 175 -1585 195
rect -1615 170 -1585 175
rect -1790 165 -1770 170
rect -1610 165 -1590 170
rect -1475 150 -1455 495
rect -1115 405 -1095 410
rect -1120 400 -1090 405
rect -1120 380 -1115 400
rect -1095 380 -1090 400
rect -1120 375 -1090 380
rect -1430 325 -1410 330
rect -1250 325 -1230 330
rect -1435 320 -1405 325
rect -1435 300 -1430 320
rect -1410 300 -1405 320
rect -1435 295 -1405 300
rect -1255 320 -1225 325
rect -1255 300 -1250 320
rect -1230 300 -1225 320
rect -1255 295 -1225 300
rect -1430 200 -1410 295
rect -1250 200 -1230 295
rect -1435 195 -1405 200
rect -1435 175 -1430 195
rect -1410 175 -1405 195
rect -1435 170 -1405 175
rect -1255 195 -1225 200
rect -1255 175 -1250 195
rect -1230 175 -1225 195
rect -1255 170 -1225 175
rect -1430 165 -1410 170
rect -1250 165 -1230 170
rect -1115 150 -1095 375
rect -1070 285 -1050 290
rect -890 285 -870 290
rect -1075 280 -1045 285
rect -1075 260 -1070 280
rect -1050 260 -1045 280
rect -1075 255 -1045 260
rect -895 280 -865 285
rect -895 260 -890 280
rect -870 260 -865 280
rect -895 255 -865 260
rect -1070 200 -1050 255
rect -890 200 -870 255
rect -1075 195 -1045 200
rect -1075 175 -1070 195
rect -1050 175 -1045 195
rect -1075 170 -1045 175
rect -895 195 -865 200
rect -895 175 -890 195
rect -870 175 -865 195
rect -895 170 -865 175
rect -1070 165 -1050 170
rect -890 165 -870 170
rect -665 150 -645 830
rect -575 725 -555 830
rect -580 720 -550 725
rect -580 700 -575 720
rect -555 700 -550 720
rect -580 695 -550 700
rect -575 150 -555 695
rect -485 565 -465 830
rect -395 645 -375 830
rect -400 640 -370 645
rect -400 620 -395 640
rect -375 620 -370 640
rect -400 615 -370 620
rect -490 560 -460 565
rect -490 540 -485 560
rect -465 540 -460 560
rect -490 535 -460 540
rect -485 150 -465 535
rect -395 150 -375 615
rect -305 605 -285 830
rect -310 600 -280 605
rect -310 580 -305 600
rect -285 580 -280 600
rect -310 575 -280 580
rect -305 150 -285 575
rect -215 325 -195 830
rect -220 320 -190 325
rect -220 300 -215 320
rect -195 300 -190 320
rect -220 295 -190 300
rect -215 150 -195 295
rect -125 285 -105 830
rect -130 280 -100 285
rect -130 260 -125 280
rect -105 260 -100 280
rect -130 255 -100 260
rect -125 150 -105 255
rect -11560 140 -11530 150
rect -11560 60 -11555 140
rect -11535 60 -11530 140
rect -11560 50 -11530 60
rect -11470 50 -11440 150
rect -11380 50 -11350 150
rect -11290 50 -11260 150
rect -11200 50 -11170 150
rect -11110 50 -11080 150
rect -11020 50 -10990 150
rect -10930 50 -10900 150
rect -10840 140 -10810 150
rect -10840 60 -10835 140
rect -10815 60 -10810 140
rect -10840 50 -10810 60
rect -10750 140 -10720 150
rect -10750 60 -10745 140
rect -10725 60 -10720 140
rect -10750 50 -10720 60
rect -10660 140 -10630 150
rect -10660 60 -10655 140
rect -10635 60 -10630 140
rect -10660 50 -10630 60
rect -10570 140 -10540 150
rect -10570 60 -10565 140
rect -10545 60 -10540 140
rect -10570 50 -10540 60
rect -10480 140 -10450 150
rect -10480 60 -10475 140
rect -10455 60 -10450 140
rect -10480 50 -10450 60
rect -10390 140 -10360 150
rect -10390 60 -10385 140
rect -10365 60 -10360 140
rect -10390 50 -10360 60
rect -10300 140 -10270 150
rect -10300 60 -10295 140
rect -10275 60 -10270 140
rect -10300 50 -10270 60
rect -10210 140 -10180 150
rect -10210 60 -10205 140
rect -10185 60 -10180 140
rect -10210 50 -10180 60
rect -10120 140 -10090 150
rect -10120 60 -10115 140
rect -10095 60 -10090 140
rect -10120 50 -10090 60
rect -10030 140 -10000 150
rect -10030 60 -10025 140
rect -10005 60 -10000 140
rect -10030 50 -10000 60
rect -9940 140 -9910 150
rect -9940 60 -9935 140
rect -9915 60 -9910 140
rect -9940 50 -9910 60
rect -9850 140 -9820 150
rect -9850 60 -9845 140
rect -9825 60 -9820 140
rect -9850 50 -9820 60
rect -9760 140 -9730 150
rect -9760 60 -9755 140
rect -9735 60 -9730 140
rect -9760 50 -9730 60
rect -9670 140 -9640 150
rect -9670 60 -9665 140
rect -9645 60 -9640 140
rect -9670 50 -9640 60
rect -9580 140 -9550 150
rect -9580 60 -9575 140
rect -9555 60 -9550 140
rect -9580 50 -9550 60
rect -9490 140 -9460 150
rect -9490 60 -9485 140
rect -9465 60 -9460 140
rect -9490 50 -9460 60
rect -9400 140 -9370 150
rect -9400 60 -9395 140
rect -9375 60 -9370 140
rect -9400 50 -9370 60
rect -9310 140 -9280 150
rect -9310 60 -9305 140
rect -9285 60 -9280 140
rect -9310 50 -9280 60
rect -9220 140 -9190 150
rect -9220 60 -9215 140
rect -9195 60 -9190 140
rect -9220 50 -9190 60
rect -9130 140 -9100 150
rect -9130 60 -9125 140
rect -9105 60 -9100 140
rect -9130 50 -9100 60
rect -9040 140 -9010 150
rect -9040 60 -9035 140
rect -9015 60 -9010 140
rect -9040 50 -9010 60
rect -8950 140 -8920 150
rect -8950 60 -8945 140
rect -8925 60 -8920 140
rect -8950 50 -8920 60
rect -8860 140 -8830 150
rect -8860 60 -8855 140
rect -8835 60 -8830 140
rect -8860 50 -8830 60
rect -8770 140 -8740 150
rect -8770 60 -8765 140
rect -8745 60 -8740 140
rect -8770 50 -8740 60
rect -8680 140 -8650 150
rect -8680 60 -8675 140
rect -8655 60 -8650 140
rect -8680 50 -8650 60
rect -8590 140 -8560 150
rect -8590 60 -8585 140
rect -8565 60 -8560 140
rect -8590 50 -8560 60
rect -8500 140 -8470 150
rect -8500 60 -8495 140
rect -8475 60 -8470 140
rect -8500 50 -8470 60
rect -8410 140 -8380 150
rect -8410 60 -8405 140
rect -8385 60 -8380 140
rect -8410 50 -8380 60
rect -8320 140 -8290 150
rect -8320 60 -8315 140
rect -8295 60 -8290 140
rect -8320 50 -8290 60
rect -8230 140 -8200 150
rect -8230 60 -8225 140
rect -8205 60 -8200 140
rect -8230 50 -8200 60
rect -8140 140 -8110 150
rect -8140 60 -8135 140
rect -8115 60 -8110 140
rect -8140 50 -8110 60
rect -8050 140 -8020 150
rect -8050 60 -8045 140
rect -8025 60 -8020 140
rect -8050 50 -8020 60
rect -7960 140 -7930 150
rect -7960 60 -7955 140
rect -7935 60 -7930 140
rect -7960 50 -7930 60
rect -7870 140 -7840 150
rect -7870 60 -7865 140
rect -7845 60 -7840 140
rect -7870 50 -7840 60
rect -7780 140 -7750 150
rect -7780 60 -7775 140
rect -7755 60 -7750 140
rect -7780 50 -7750 60
rect -7690 140 -7660 150
rect -7690 60 -7685 140
rect -7665 60 -7660 140
rect -7690 50 -7660 60
rect -7600 140 -7570 150
rect -7600 60 -7595 140
rect -7575 60 -7570 140
rect -7600 50 -7570 60
rect -7510 140 -7480 150
rect -7510 60 -7505 140
rect -7485 60 -7480 140
rect -7510 50 -7480 60
rect -7420 140 -7390 150
rect -7420 60 -7415 140
rect -7395 60 -7390 140
rect -7420 50 -7390 60
rect -7330 140 -7300 150
rect -7330 60 -7325 140
rect -7305 60 -7300 140
rect -7330 50 -7300 60
rect -7240 140 -7210 150
rect -7240 60 -7235 140
rect -7215 60 -7210 140
rect -7240 50 -7210 60
rect -7150 140 -7120 150
rect -7150 60 -7145 140
rect -7125 60 -7120 140
rect -7150 50 -7120 60
rect -7060 140 -7030 150
rect -7060 60 -7055 140
rect -7035 60 -7030 140
rect -7060 50 -7030 60
rect -6970 140 -6940 150
rect -6970 60 -6965 140
rect -6945 60 -6940 140
rect -6970 50 -6940 60
rect -6880 140 -6850 150
rect -6880 60 -6875 140
rect -6855 60 -6850 140
rect -6880 50 -6850 60
rect -6790 140 -6760 150
rect -6790 60 -6785 140
rect -6765 60 -6760 140
rect -6790 50 -6760 60
rect -6700 140 -6670 150
rect -6700 60 -6695 140
rect -6675 60 -6670 140
rect -6700 50 -6670 60
rect -6610 140 -6580 150
rect -6610 60 -6605 140
rect -6585 60 -6580 140
rect -6610 50 -6580 60
rect -6520 140 -6490 150
rect -6520 60 -6515 140
rect -6495 60 -6490 140
rect -6520 50 -6490 60
rect -6430 140 -6400 150
rect -6430 60 -6425 140
rect -6405 60 -6400 140
rect -6430 50 -6400 60
rect -6340 140 -6310 150
rect -6340 60 -6335 140
rect -6315 60 -6310 140
rect -6340 50 -6310 60
rect -6250 140 -6220 150
rect -6250 60 -6245 140
rect -6225 60 -6220 140
rect -6250 50 -6220 60
rect -6160 140 -6130 150
rect -6160 60 -6155 140
rect -6135 60 -6130 140
rect -6160 50 -6130 60
rect -6070 140 -6040 150
rect -6070 60 -6065 140
rect -6045 60 -6040 140
rect -6070 50 -6040 60
rect -5980 140 -5950 150
rect -5980 60 -5975 140
rect -5955 60 -5950 140
rect -5980 50 -5950 60
rect -5890 140 -5860 150
rect -5890 60 -5885 140
rect -5865 60 -5860 140
rect -5890 50 -5860 60
rect -5800 140 -5770 150
rect -5800 60 -5795 140
rect -5775 60 -5770 140
rect -5800 50 -5770 60
rect -5710 140 -5680 150
rect -5710 60 -5705 140
rect -5685 60 -5680 140
rect -5710 50 -5680 60
rect -5620 140 -5590 150
rect -5620 60 -5615 140
rect -5595 60 -5590 140
rect -5620 50 -5590 60
rect -5530 140 -5500 150
rect -5530 60 -5525 140
rect -5505 60 -5500 140
rect -5530 50 -5500 60
rect -5440 140 -5410 150
rect -5440 60 -5435 140
rect -5415 60 -5410 140
rect -5440 50 -5410 60
rect -5350 140 -5320 150
rect -5350 60 -5345 140
rect -5325 60 -5320 140
rect -5350 50 -5320 60
rect -5260 140 -5230 150
rect -5260 60 -5255 140
rect -5235 60 -5230 140
rect -5260 50 -5230 60
rect -5170 140 -5140 150
rect -5170 60 -5165 140
rect -5145 60 -5140 140
rect -5170 50 -5140 60
rect -5080 140 -5050 150
rect -5080 60 -5075 140
rect -5055 60 -5050 140
rect -5080 50 -5050 60
rect -4990 140 -4960 150
rect -4990 60 -4985 140
rect -4965 60 -4960 140
rect -4990 50 -4960 60
rect -4900 140 -4870 150
rect -4900 60 -4895 140
rect -4875 60 -4870 140
rect -4900 50 -4870 60
rect -4810 140 -4780 150
rect -4810 60 -4805 140
rect -4785 60 -4780 140
rect -4810 50 -4780 60
rect -4720 140 -4690 150
rect -4720 60 -4715 140
rect -4695 60 -4690 140
rect -4720 50 -4690 60
rect -4630 140 -4600 150
rect -4630 60 -4625 140
rect -4605 60 -4600 140
rect -4630 50 -4600 60
rect -4540 140 -4510 150
rect -4540 60 -4535 140
rect -4515 60 -4510 140
rect -4540 50 -4510 60
rect -4450 140 -4420 150
rect -4450 60 -4445 140
rect -4425 60 -4420 140
rect -4450 50 -4420 60
rect -4360 140 -4330 150
rect -4360 60 -4355 140
rect -4335 60 -4330 140
rect -4360 50 -4330 60
rect -4270 140 -4240 150
rect -4270 60 -4265 140
rect -4245 60 -4240 140
rect -4270 50 -4240 60
rect -4180 140 -4150 150
rect -4180 60 -4175 140
rect -4155 60 -4150 140
rect -4180 50 -4150 60
rect -4090 140 -4060 150
rect -4090 60 -4085 140
rect -4065 60 -4060 140
rect -4090 50 -4060 60
rect -4000 140 -3970 150
rect -4000 60 -3995 140
rect -3975 60 -3970 140
rect -4000 50 -3970 60
rect -3910 140 -3880 150
rect -3910 60 -3905 140
rect -3885 60 -3880 140
rect -3910 50 -3880 60
rect -3820 140 -3790 150
rect -3820 60 -3815 140
rect -3795 60 -3790 140
rect -3820 50 -3790 60
rect -3730 140 -3700 150
rect -3730 60 -3725 140
rect -3705 60 -3700 140
rect -3730 50 -3700 60
rect -3640 140 -3610 150
rect -3640 60 -3635 140
rect -3615 60 -3610 140
rect -3640 50 -3610 60
rect -3550 140 -3520 150
rect -3550 60 -3545 140
rect -3525 60 -3520 140
rect -3550 50 -3520 60
rect -3460 140 -3430 150
rect -3460 60 -3455 140
rect -3435 60 -3430 140
rect -3460 50 -3430 60
rect -3370 140 -3340 150
rect -3370 60 -3365 140
rect -3345 60 -3340 140
rect -3370 50 -3340 60
rect -3280 140 -3250 150
rect -3280 60 -3275 140
rect -3255 60 -3250 140
rect -3280 50 -3250 60
rect -3190 140 -3160 150
rect -3190 60 -3185 140
rect -3165 60 -3160 140
rect -3190 50 -3160 60
rect -3100 140 -3070 150
rect -3100 60 -3095 140
rect -3075 60 -3070 140
rect -3100 50 -3070 60
rect -3010 140 -2980 150
rect -3010 60 -3005 140
rect -2985 60 -2980 140
rect -3010 50 -2980 60
rect -2920 140 -2890 150
rect -2920 60 -2915 140
rect -2895 60 -2890 140
rect -2920 50 -2890 60
rect -2830 140 -2800 150
rect -2830 60 -2825 140
rect -2805 60 -2800 140
rect -2830 50 -2800 60
rect -2740 140 -2710 150
rect -2740 60 -2735 140
rect -2715 60 -2710 140
rect -2740 50 -2710 60
rect -2650 140 -2620 150
rect -2650 60 -2645 140
rect -2625 60 -2620 140
rect -2650 50 -2620 60
rect -2560 140 -2530 150
rect -2560 60 -2555 140
rect -2535 60 -2530 140
rect -2560 50 -2530 60
rect -2470 140 -2440 150
rect -2470 60 -2465 140
rect -2445 60 -2440 140
rect -2470 50 -2440 60
rect -2380 140 -2350 150
rect -2380 60 -2375 140
rect -2355 60 -2350 140
rect -2380 50 -2350 60
rect -2290 140 -2260 150
rect -2290 60 -2285 140
rect -2265 60 -2260 140
rect -2290 50 -2260 60
rect -2200 140 -2170 150
rect -2200 60 -2195 140
rect -2175 60 -2170 140
rect -2200 50 -2170 60
rect -2110 140 -2080 150
rect -2110 60 -2105 140
rect -2085 60 -2080 140
rect -2110 50 -2080 60
rect -2020 140 -1990 150
rect -2020 60 -2015 140
rect -1995 60 -1990 140
rect -2020 50 -1990 60
rect -1930 140 -1900 150
rect -1930 60 -1925 140
rect -1905 60 -1900 140
rect -1930 50 -1900 60
rect -1840 140 -1810 150
rect -1840 60 -1835 140
rect -1815 60 -1810 140
rect -1840 50 -1810 60
rect -1750 140 -1720 150
rect -1750 60 -1745 140
rect -1725 60 -1720 140
rect -1750 50 -1720 60
rect -1660 140 -1630 150
rect -1660 60 -1655 140
rect -1635 60 -1630 140
rect -1660 50 -1630 60
rect -1570 140 -1540 150
rect -1570 60 -1565 140
rect -1545 60 -1540 140
rect -1570 50 -1540 60
rect -1480 140 -1450 150
rect -1480 60 -1475 140
rect -1455 60 -1450 140
rect -1480 50 -1450 60
rect -1390 140 -1360 150
rect -1390 60 -1385 140
rect -1365 60 -1360 140
rect -1390 50 -1360 60
rect -1300 140 -1270 150
rect -1300 60 -1295 140
rect -1275 60 -1270 140
rect -1300 50 -1270 60
rect -1210 140 -1180 150
rect -1210 60 -1205 140
rect -1185 60 -1180 140
rect -1210 50 -1180 60
rect -1120 140 -1090 150
rect -1120 60 -1115 140
rect -1095 60 -1090 140
rect -1120 50 -1090 60
rect -1030 140 -1000 150
rect -1030 60 -1025 140
rect -1005 60 -1000 140
rect -1030 50 -1000 60
rect -940 140 -910 150
rect -940 60 -935 140
rect -915 60 -910 140
rect -940 50 -910 60
rect -850 140 -820 150
rect -850 60 -845 140
rect -825 60 -820 140
rect -850 50 -820 60
rect -760 140 -730 150
rect -760 60 -755 140
rect -735 60 -730 140
rect -760 50 -730 60
rect -670 50 -640 150
rect -580 50 -550 150
rect -490 50 -460 150
rect -400 50 -370 150
rect -310 50 -280 150
rect -220 50 -190 150
rect -130 50 -100 150
rect -40 140 -10 150
rect -40 60 -35 140
rect -15 60 -10 140
rect -40 50 -10 60
rect -11555 30 -11535 50
rect -10835 30 -10815 50
rect -7235 30 -7215 50
rect -3635 30 -3615 50
rect -2195 30 -2175 50
rect -755 30 -735 50
rect -35 30 -15 50
rect -11700 -5 -11695 25
rect -11665 -5 -11660 25
rect -11700 -10 -11660 -5
rect -11565 25 -11525 30
rect -11565 -5 -11560 25
rect -11530 -5 -11525 25
rect -11565 -10 -11525 -5
rect -10845 25 -10805 30
rect -10845 -5 -10840 25
rect -10810 -5 -10805 25
rect -10845 -10 -10805 -5
rect -10665 25 -10625 30
rect -10665 -5 -10660 25
rect -10630 -5 -10625 25
rect -10665 -10 -10625 -5
rect -10485 25 -10445 30
rect -10485 -5 -10480 25
rect -10450 -5 -10445 25
rect -10485 -10 -10445 -5
rect -10305 25 -10265 30
rect -10305 -5 -10300 25
rect -10270 -5 -10265 25
rect -10305 -10 -10265 -5
rect -10125 25 -10085 30
rect -10125 -5 -10120 25
rect -10090 -5 -10085 25
rect -10125 -10 -10085 -5
rect -9945 25 -9905 30
rect -9945 -5 -9940 25
rect -9910 -5 -9905 25
rect -9945 -10 -9905 -5
rect -9765 25 -9725 30
rect -9765 -5 -9760 25
rect -9730 -5 -9725 25
rect -9765 -10 -9725 -5
rect -9585 25 -9545 30
rect -9585 -5 -9580 25
rect -9550 -5 -9545 25
rect -9585 -10 -9545 -5
rect -9405 25 -9365 30
rect -9405 -5 -9400 25
rect -9370 -5 -9365 25
rect -9405 -10 -9365 -5
rect -9225 25 -9185 30
rect -9225 -5 -9220 25
rect -9190 -5 -9185 25
rect -9225 -10 -9185 -5
rect -9045 25 -9005 30
rect -9045 -5 -9040 25
rect -9010 -5 -9005 25
rect -9045 -10 -9005 -5
rect -8865 25 -8825 30
rect -8865 -5 -8860 25
rect -8830 -5 -8825 25
rect -8865 -10 -8825 -5
rect -8685 25 -8645 30
rect -8685 -5 -8680 25
rect -8650 -5 -8645 25
rect -8685 -10 -8645 -5
rect -8505 25 -8465 30
rect -8505 -5 -8500 25
rect -8470 -5 -8465 25
rect -8505 -10 -8465 -5
rect -8325 25 -8285 30
rect -8325 -5 -8320 25
rect -8290 -5 -8285 25
rect -8325 -10 -8285 -5
rect -8145 25 -8105 30
rect -8145 -5 -8140 25
rect -8110 -5 -8105 25
rect -8145 -10 -8105 -5
rect -7965 25 -7925 30
rect -7965 -5 -7960 25
rect -7930 -5 -7925 25
rect -7965 -10 -7925 -5
rect -7785 25 -7745 30
rect -7785 -5 -7780 25
rect -7750 -5 -7745 25
rect -7785 -10 -7745 -5
rect -7605 25 -7565 30
rect -7605 -5 -7600 25
rect -7570 -5 -7565 25
rect -7605 -10 -7565 -5
rect -7425 25 -7385 30
rect -7425 -5 -7420 25
rect -7390 -5 -7385 25
rect -7425 -10 -7385 -5
rect -7245 25 -7205 30
rect -7245 -5 -7240 25
rect -7210 -5 -7205 25
rect -7245 -10 -7205 -5
rect -7065 25 -7025 30
rect -7065 -5 -7060 25
rect -7030 -5 -7025 25
rect -7065 -10 -7025 -5
rect -6885 25 -6845 30
rect -6885 -5 -6880 25
rect -6850 -5 -6845 25
rect -6885 -10 -6845 -5
rect -6705 25 -6665 30
rect -6705 -5 -6700 25
rect -6670 -5 -6665 25
rect -6705 -10 -6665 -5
rect -6525 25 -6485 30
rect -6525 -5 -6520 25
rect -6490 -5 -6485 25
rect -6525 -10 -6485 -5
rect -6345 25 -6305 30
rect -6345 -5 -6340 25
rect -6310 -5 -6305 25
rect -6345 -10 -6305 -5
rect -6165 25 -6125 30
rect -6165 -5 -6160 25
rect -6130 -5 -6125 25
rect -6165 -10 -6125 -5
rect -5985 25 -5945 30
rect -5985 -5 -5980 25
rect -5950 -5 -5945 25
rect -5985 -10 -5945 -5
rect -5805 25 -5765 30
rect -5805 -5 -5800 25
rect -5770 -5 -5765 25
rect -5805 -10 -5765 -5
rect -5625 25 -5585 30
rect -5625 -5 -5620 25
rect -5590 -5 -5585 25
rect -5625 -10 -5585 -5
rect -5445 25 -5405 30
rect -5445 -5 -5440 25
rect -5410 -5 -5405 25
rect -5445 -10 -5405 -5
rect -5265 25 -5225 30
rect -5265 -5 -5260 25
rect -5230 -5 -5225 25
rect -5265 -10 -5225 -5
rect -5085 25 -5045 30
rect -5085 -5 -5080 25
rect -5050 -5 -5045 25
rect -5085 -10 -5045 -5
rect -4905 25 -4865 30
rect -4905 -5 -4900 25
rect -4870 -5 -4865 25
rect -4905 -10 -4865 -5
rect -4725 25 -4685 30
rect -4725 -5 -4720 25
rect -4690 -5 -4685 25
rect -4725 -10 -4685 -5
rect -4545 25 -4505 30
rect -4545 -5 -4540 25
rect -4510 -5 -4505 25
rect -4545 -10 -4505 -5
rect -4365 25 -4325 30
rect -4365 -5 -4360 25
rect -4330 -5 -4325 25
rect -4365 -10 -4325 -5
rect -4185 25 -4145 30
rect -4185 -5 -4180 25
rect -4150 -5 -4145 25
rect -4185 -10 -4145 -5
rect -4005 25 -3965 30
rect -4005 -5 -4000 25
rect -3970 -5 -3965 25
rect -4005 -10 -3965 -5
rect -3825 25 -3785 30
rect -3825 -5 -3820 25
rect -3790 -5 -3785 25
rect -3825 -10 -3785 -5
rect -3645 25 -3605 30
rect -3645 -5 -3640 25
rect -3610 -5 -3605 25
rect -3645 -10 -3605 -5
rect -3465 25 -3425 30
rect -3465 -5 -3460 25
rect -3430 -5 -3425 25
rect -3465 -10 -3425 -5
rect -3285 25 -3245 30
rect -3285 -5 -3280 25
rect -3250 -5 -3245 25
rect -3285 -10 -3245 -5
rect -3105 25 -3065 30
rect -3105 -5 -3100 25
rect -3070 -5 -3065 25
rect -3105 -10 -3065 -5
rect -2925 25 -2885 30
rect -2925 -5 -2920 25
rect -2890 -5 -2885 25
rect -2925 -10 -2885 -5
rect -2745 25 -2705 30
rect -2745 -5 -2740 25
rect -2710 -5 -2705 25
rect -2745 -10 -2705 -5
rect -2565 25 -2525 30
rect -2565 -5 -2560 25
rect -2530 -5 -2525 25
rect -2565 -10 -2525 -5
rect -2385 25 -2345 30
rect -2385 -5 -2380 25
rect -2350 -5 -2345 25
rect -2385 -10 -2345 -5
rect -2205 25 -2165 30
rect -2205 -5 -2200 25
rect -2170 -5 -2165 25
rect -2205 -10 -2165 -5
rect -2025 25 -1985 30
rect -2025 -5 -2020 25
rect -1990 -5 -1985 25
rect -2025 -10 -1985 -5
rect -1845 25 -1805 30
rect -1845 -5 -1840 25
rect -1810 -5 -1805 25
rect -1845 -10 -1805 -5
rect -1665 25 -1625 30
rect -1665 -5 -1660 25
rect -1630 -5 -1625 25
rect -1665 -10 -1625 -5
rect -1485 25 -1445 30
rect -1485 -5 -1480 25
rect -1450 -5 -1445 25
rect -1485 -10 -1445 -5
rect -1305 25 -1265 30
rect -1305 -5 -1300 25
rect -1270 -5 -1265 25
rect -1305 -10 -1265 -5
rect -1125 25 -1085 30
rect -1125 -5 -1120 25
rect -1090 -5 -1085 25
rect -1125 -10 -1085 -5
rect -945 25 -905 30
rect -945 -5 -940 25
rect -910 -5 -905 25
rect -945 -10 -905 -5
rect -765 25 -725 30
rect -765 -5 -760 25
rect -730 -5 -725 25
rect -765 -10 -725 -5
rect -45 25 -5 30
rect -45 -5 -40 25
rect -10 -5 -5 25
rect -45 -10 -5 -5
rect 90 25 130 1970
rect 90 -5 95 25
rect 125 -5 130 25
rect 90 -10 130 -5
<< via1 >>
rect -11695 1995 -11665 2000
rect -11695 1975 -11690 1995
rect -11690 1975 -11670 1995
rect -11670 1975 -11665 1995
rect -11695 1970 -11665 1975
rect -11560 1995 -11530 2000
rect -11560 1975 -11555 1995
rect -11555 1975 -11535 1995
rect -11535 1975 -11530 1995
rect -11560 1970 -11530 1975
rect -10840 1995 -10810 2000
rect -10840 1975 -10835 1995
rect -10835 1975 -10815 1995
rect -10815 1975 -10810 1995
rect -10840 1970 -10810 1975
rect -10660 1995 -10630 2000
rect -10660 1975 -10655 1995
rect -10655 1975 -10635 1995
rect -10635 1975 -10630 1995
rect -10660 1970 -10630 1975
rect -10480 1995 -10450 2000
rect -10480 1975 -10475 1995
rect -10475 1975 -10455 1995
rect -10455 1975 -10450 1995
rect -10480 1970 -10450 1975
rect -10300 1995 -10270 2000
rect -10300 1975 -10295 1995
rect -10295 1975 -10275 1995
rect -10275 1975 -10270 1995
rect -10300 1970 -10270 1975
rect -10120 1995 -10090 2000
rect -10120 1975 -10115 1995
rect -10115 1975 -10095 1995
rect -10095 1975 -10090 1995
rect -10120 1970 -10090 1975
rect -9940 1995 -9910 2000
rect -9940 1975 -9935 1995
rect -9935 1975 -9915 1995
rect -9915 1975 -9910 1995
rect -9940 1970 -9910 1975
rect -9760 1995 -9730 2000
rect -9760 1975 -9755 1995
rect -9755 1975 -9735 1995
rect -9735 1975 -9730 1995
rect -9760 1970 -9730 1975
rect -9580 1995 -9550 2000
rect -9580 1975 -9575 1995
rect -9575 1975 -9555 1995
rect -9555 1975 -9550 1995
rect -9580 1970 -9550 1975
rect -9400 1995 -9370 2000
rect -9400 1975 -9395 1995
rect -9395 1975 -9375 1995
rect -9375 1975 -9370 1995
rect -9400 1970 -9370 1975
rect -9220 1995 -9190 2000
rect -9220 1975 -9215 1995
rect -9215 1975 -9195 1995
rect -9195 1975 -9190 1995
rect -9220 1970 -9190 1975
rect -9040 1995 -9010 2000
rect -9040 1975 -9035 1995
rect -9035 1975 -9015 1995
rect -9015 1975 -9010 1995
rect -9040 1970 -9010 1975
rect -8860 1995 -8830 2000
rect -8860 1975 -8855 1995
rect -8855 1975 -8835 1995
rect -8835 1975 -8830 1995
rect -8860 1970 -8830 1975
rect -8680 1995 -8650 2000
rect -8680 1975 -8675 1995
rect -8675 1975 -8655 1995
rect -8655 1975 -8650 1995
rect -8680 1970 -8650 1975
rect -8500 1995 -8470 2000
rect -8500 1975 -8495 1995
rect -8495 1975 -8475 1995
rect -8475 1975 -8470 1995
rect -8500 1970 -8470 1975
rect -8320 1995 -8290 2000
rect -8320 1975 -8315 1995
rect -8315 1975 -8295 1995
rect -8295 1975 -8290 1995
rect -8320 1970 -8290 1975
rect -8140 1995 -8110 2000
rect -8140 1975 -8135 1995
rect -8135 1975 -8115 1995
rect -8115 1975 -8110 1995
rect -8140 1970 -8110 1975
rect -7960 1995 -7930 2000
rect -7960 1975 -7955 1995
rect -7955 1975 -7935 1995
rect -7935 1975 -7930 1995
rect -7960 1970 -7930 1975
rect -7780 1995 -7750 2000
rect -7780 1975 -7775 1995
rect -7775 1975 -7755 1995
rect -7755 1975 -7750 1995
rect -7780 1970 -7750 1975
rect -7600 1995 -7570 2000
rect -7600 1975 -7595 1995
rect -7595 1975 -7575 1995
rect -7575 1975 -7570 1995
rect -7600 1970 -7570 1975
rect -7420 1995 -7390 2000
rect -7420 1975 -7415 1995
rect -7415 1975 -7395 1995
rect -7395 1975 -7390 1995
rect -7420 1970 -7390 1975
rect -7240 1995 -7210 2000
rect -7240 1975 -7235 1995
rect -7235 1975 -7215 1995
rect -7215 1975 -7210 1995
rect -7240 1970 -7210 1975
rect -7060 1995 -7030 2000
rect -7060 1975 -7055 1995
rect -7055 1975 -7035 1995
rect -7035 1975 -7030 1995
rect -7060 1970 -7030 1975
rect -6880 1995 -6850 2000
rect -6880 1975 -6875 1995
rect -6875 1975 -6855 1995
rect -6855 1975 -6850 1995
rect -6880 1970 -6850 1975
rect -6700 1995 -6670 2000
rect -6700 1975 -6695 1995
rect -6695 1975 -6675 1995
rect -6675 1975 -6670 1995
rect -6700 1970 -6670 1975
rect -6520 1995 -6490 2000
rect -6520 1975 -6515 1995
rect -6515 1975 -6495 1995
rect -6495 1975 -6490 1995
rect -6520 1970 -6490 1975
rect -6340 1995 -6310 2000
rect -6340 1975 -6335 1995
rect -6335 1975 -6315 1995
rect -6315 1975 -6310 1995
rect -6340 1970 -6310 1975
rect -6160 1995 -6130 2000
rect -6160 1975 -6155 1995
rect -6155 1975 -6135 1995
rect -6135 1975 -6130 1995
rect -6160 1970 -6130 1975
rect -5980 1995 -5950 2000
rect -5980 1975 -5975 1995
rect -5975 1975 -5955 1995
rect -5955 1975 -5950 1995
rect -5980 1970 -5950 1975
rect -5800 1995 -5770 2000
rect -5800 1975 -5795 1995
rect -5795 1975 -5775 1995
rect -5775 1975 -5770 1995
rect -5800 1970 -5770 1975
rect -5620 1995 -5590 2000
rect -5620 1975 -5615 1995
rect -5615 1975 -5595 1995
rect -5595 1975 -5590 1995
rect -5620 1970 -5590 1975
rect -5440 1995 -5410 2000
rect -5440 1975 -5435 1995
rect -5435 1975 -5415 1995
rect -5415 1975 -5410 1995
rect -5440 1970 -5410 1975
rect -5260 1995 -5230 2000
rect -5260 1975 -5255 1995
rect -5255 1975 -5235 1995
rect -5235 1975 -5230 1995
rect -5260 1970 -5230 1975
rect -5080 1995 -5050 2000
rect -5080 1975 -5075 1995
rect -5075 1975 -5055 1995
rect -5055 1975 -5050 1995
rect -5080 1970 -5050 1975
rect -4900 1995 -4870 2000
rect -4900 1975 -4895 1995
rect -4895 1975 -4875 1995
rect -4875 1975 -4870 1995
rect -4900 1970 -4870 1975
rect -4720 1995 -4690 2000
rect -4720 1975 -4715 1995
rect -4715 1975 -4695 1995
rect -4695 1975 -4690 1995
rect -4720 1970 -4690 1975
rect -4540 1995 -4510 2000
rect -4540 1975 -4535 1995
rect -4535 1975 -4515 1995
rect -4515 1975 -4510 1995
rect -4540 1970 -4510 1975
rect -4360 1995 -4330 2000
rect -4360 1975 -4355 1995
rect -4355 1975 -4335 1995
rect -4335 1975 -4330 1995
rect -4360 1970 -4330 1975
rect -4180 1995 -4150 2000
rect -4180 1975 -4175 1995
rect -4175 1975 -4155 1995
rect -4155 1975 -4150 1995
rect -4180 1970 -4150 1975
rect -4000 1995 -3970 2000
rect -4000 1975 -3995 1995
rect -3995 1975 -3975 1995
rect -3975 1975 -3970 1995
rect -4000 1970 -3970 1975
rect -3820 1995 -3790 2000
rect -3820 1975 -3815 1995
rect -3815 1975 -3795 1995
rect -3795 1975 -3790 1995
rect -3820 1970 -3790 1975
rect -3640 1995 -3610 2000
rect -3640 1975 -3635 1995
rect -3635 1975 -3615 1995
rect -3615 1975 -3610 1995
rect -3640 1970 -3610 1975
rect -3460 1995 -3430 2000
rect -3460 1975 -3455 1995
rect -3455 1975 -3435 1995
rect -3435 1975 -3430 1995
rect -3460 1970 -3430 1975
rect -3280 1995 -3250 2000
rect -3280 1975 -3275 1995
rect -3275 1975 -3255 1995
rect -3255 1975 -3250 1995
rect -3280 1970 -3250 1975
rect -3100 1995 -3070 2000
rect -3100 1975 -3095 1995
rect -3095 1975 -3075 1995
rect -3075 1975 -3070 1995
rect -3100 1970 -3070 1975
rect -2920 1995 -2890 2000
rect -2920 1975 -2915 1995
rect -2915 1975 -2895 1995
rect -2895 1975 -2890 1995
rect -2920 1970 -2890 1975
rect -2740 1995 -2710 2000
rect -2740 1975 -2735 1995
rect -2735 1975 -2715 1995
rect -2715 1975 -2710 1995
rect -2740 1970 -2710 1975
rect -2560 1995 -2530 2000
rect -2560 1975 -2555 1995
rect -2555 1975 -2535 1995
rect -2535 1975 -2530 1995
rect -2560 1970 -2530 1975
rect -2380 1995 -2350 2000
rect -2380 1975 -2375 1995
rect -2375 1975 -2355 1995
rect -2355 1975 -2350 1995
rect -2380 1970 -2350 1975
rect -2200 1995 -2170 2000
rect -2200 1975 -2195 1995
rect -2195 1975 -2175 1995
rect -2175 1975 -2170 1995
rect -2200 1970 -2170 1975
rect -2020 1995 -1990 2000
rect -2020 1975 -2015 1995
rect -2015 1975 -1995 1995
rect -1995 1975 -1990 1995
rect -2020 1970 -1990 1975
rect -1840 1995 -1810 2000
rect -1840 1975 -1835 1995
rect -1835 1975 -1815 1995
rect -1815 1975 -1810 1995
rect -1840 1970 -1810 1975
rect -1660 1995 -1630 2000
rect -1660 1975 -1655 1995
rect -1655 1975 -1635 1995
rect -1635 1975 -1630 1995
rect -1660 1970 -1630 1975
rect -1480 1995 -1450 2000
rect -1480 1975 -1475 1995
rect -1475 1975 -1455 1995
rect -1455 1975 -1450 1995
rect -1480 1970 -1450 1975
rect -1300 1995 -1270 2000
rect -1300 1975 -1295 1995
rect -1295 1975 -1275 1995
rect -1275 1975 -1270 1995
rect -1300 1970 -1270 1975
rect -1120 1995 -1090 2000
rect -1120 1975 -1115 1995
rect -1115 1975 -1095 1995
rect -1095 1975 -1090 1995
rect -1120 1970 -1090 1975
rect -940 1995 -910 2000
rect -940 1975 -935 1995
rect -935 1975 -915 1995
rect -915 1975 -910 1995
rect -940 1970 -910 1975
rect -760 1995 -730 2000
rect -760 1975 -755 1995
rect -755 1975 -735 1995
rect -735 1975 -730 1995
rect -760 1970 -730 1975
rect -40 1995 -10 2000
rect -40 1975 -35 1995
rect -35 1975 -15 1995
rect -15 1975 -10 1995
rect -40 1970 -10 1975
rect 95 1995 125 2000
rect 95 1975 100 1995
rect 100 1975 120 1995
rect 120 1975 125 1995
rect 95 1970 125 1975
rect -11560 1035 -11530 1040
rect -11560 1015 -11555 1035
rect -11555 1015 -11535 1035
rect -11535 1015 -11530 1035
rect -11560 1010 -11530 1015
rect -11560 980 -11530 985
rect -11560 960 -11555 980
rect -11555 960 -11535 980
rect -11535 960 -11530 980
rect -11560 955 -11530 960
rect -10840 1035 -10810 1040
rect -10840 1015 -10835 1035
rect -10835 1015 -10815 1035
rect -10815 1015 -10810 1035
rect -10840 1010 -10810 1015
rect -10660 1035 -10630 1040
rect -10660 1015 -10655 1035
rect -10655 1015 -10635 1035
rect -10635 1015 -10630 1035
rect -10660 1010 -10630 1015
rect -10480 1035 -10450 1040
rect -10480 1015 -10475 1035
rect -10475 1015 -10455 1035
rect -10455 1015 -10450 1035
rect -10480 1010 -10450 1015
rect -10300 1035 -10270 1040
rect -10300 1015 -10295 1035
rect -10295 1015 -10275 1035
rect -10275 1015 -10270 1035
rect -10300 1010 -10270 1015
rect -10120 1035 -10090 1040
rect -10120 1015 -10115 1035
rect -10115 1015 -10095 1035
rect -10095 1015 -10090 1035
rect -10120 1010 -10090 1015
rect -9940 1035 -9910 1040
rect -9940 1015 -9935 1035
rect -9935 1015 -9915 1035
rect -9915 1015 -9910 1035
rect -9940 1010 -9910 1015
rect -9760 1035 -9730 1040
rect -9760 1015 -9755 1035
rect -9755 1015 -9735 1035
rect -9735 1015 -9730 1035
rect -9760 1010 -9730 1015
rect -9580 1035 -9550 1040
rect -9580 1015 -9575 1035
rect -9575 1015 -9555 1035
rect -9555 1015 -9550 1035
rect -9580 1010 -9550 1015
rect -9400 1035 -9370 1040
rect -9400 1015 -9395 1035
rect -9395 1015 -9375 1035
rect -9375 1015 -9370 1035
rect -9400 1010 -9370 1015
rect -9220 1035 -9190 1040
rect -9220 1015 -9215 1035
rect -9215 1015 -9195 1035
rect -9195 1015 -9190 1035
rect -9220 1010 -9190 1015
rect -9040 1035 -9010 1040
rect -9040 1015 -9035 1035
rect -9035 1015 -9015 1035
rect -9015 1015 -9010 1035
rect -9040 1010 -9010 1015
rect -8860 1035 -8830 1040
rect -8860 1015 -8855 1035
rect -8855 1015 -8835 1035
rect -8835 1015 -8830 1035
rect -8860 1010 -8830 1015
rect -8680 1035 -8650 1040
rect -8680 1015 -8675 1035
rect -8675 1015 -8655 1035
rect -8655 1015 -8650 1035
rect -8680 1010 -8650 1015
rect -8500 1035 -8470 1040
rect -8500 1015 -8495 1035
rect -8495 1015 -8475 1035
rect -8475 1015 -8470 1035
rect -8500 1010 -8470 1015
rect -8320 1035 -8290 1040
rect -8320 1015 -8315 1035
rect -8315 1015 -8295 1035
rect -8295 1015 -8290 1035
rect -8320 1010 -8290 1015
rect -8140 1035 -8110 1040
rect -8140 1015 -8135 1035
rect -8135 1015 -8115 1035
rect -8115 1015 -8110 1035
rect -8140 1010 -8110 1015
rect -7960 1035 -7930 1040
rect -7960 1015 -7955 1035
rect -7955 1015 -7935 1035
rect -7935 1015 -7930 1035
rect -7960 1010 -7930 1015
rect -7780 1035 -7750 1040
rect -7780 1015 -7775 1035
rect -7775 1015 -7755 1035
rect -7755 1015 -7750 1035
rect -7780 1010 -7750 1015
rect -7600 1035 -7570 1040
rect -7600 1015 -7595 1035
rect -7595 1015 -7575 1035
rect -7575 1015 -7570 1035
rect -7600 1010 -7570 1015
rect -7420 1035 -7390 1040
rect -7420 1015 -7415 1035
rect -7415 1015 -7395 1035
rect -7395 1015 -7390 1035
rect -7420 1010 -7390 1015
rect -7240 1035 -7210 1040
rect -7240 1015 -7235 1035
rect -7235 1015 -7215 1035
rect -7215 1015 -7210 1035
rect -7240 1010 -7210 1015
rect -7060 1035 -7030 1040
rect -7060 1015 -7055 1035
rect -7055 1015 -7035 1035
rect -7035 1015 -7030 1035
rect -7060 1010 -7030 1015
rect -6880 1035 -6850 1040
rect -6880 1015 -6875 1035
rect -6875 1015 -6855 1035
rect -6855 1015 -6850 1035
rect -6880 1010 -6850 1015
rect -6700 1035 -6670 1040
rect -6700 1015 -6695 1035
rect -6695 1015 -6675 1035
rect -6675 1015 -6670 1035
rect -6700 1010 -6670 1015
rect -6520 1035 -6490 1040
rect -6520 1015 -6515 1035
rect -6515 1015 -6495 1035
rect -6495 1015 -6490 1035
rect -6520 1010 -6490 1015
rect -6340 1035 -6310 1040
rect -6340 1015 -6335 1035
rect -6335 1015 -6315 1035
rect -6315 1015 -6310 1035
rect -6340 1010 -6310 1015
rect -6160 1035 -6130 1040
rect -6160 1015 -6155 1035
rect -6155 1015 -6135 1035
rect -6135 1015 -6130 1035
rect -6160 1010 -6130 1015
rect -5980 1035 -5950 1040
rect -5980 1015 -5975 1035
rect -5975 1015 -5955 1035
rect -5955 1015 -5950 1035
rect -5980 1010 -5950 1015
rect -5800 1035 -5770 1040
rect -5800 1015 -5795 1035
rect -5795 1015 -5775 1035
rect -5775 1015 -5770 1035
rect -5800 1010 -5770 1015
rect -5620 1035 -5590 1040
rect -5620 1015 -5615 1035
rect -5615 1015 -5595 1035
rect -5595 1015 -5590 1035
rect -5620 1010 -5590 1015
rect -5440 1035 -5410 1040
rect -5440 1015 -5435 1035
rect -5435 1015 -5415 1035
rect -5415 1015 -5410 1035
rect -5440 1010 -5410 1015
rect -5260 1035 -5230 1040
rect -5260 1015 -5255 1035
rect -5255 1015 -5235 1035
rect -5235 1015 -5230 1035
rect -5260 1010 -5230 1015
rect -5080 1035 -5050 1040
rect -5080 1015 -5075 1035
rect -5075 1015 -5055 1035
rect -5055 1015 -5050 1035
rect -5080 1010 -5050 1015
rect -4900 1035 -4870 1040
rect -4900 1015 -4895 1035
rect -4895 1015 -4875 1035
rect -4875 1015 -4870 1035
rect -4900 1010 -4870 1015
rect -4720 1035 -4690 1040
rect -4720 1015 -4715 1035
rect -4715 1015 -4695 1035
rect -4695 1015 -4690 1035
rect -4720 1010 -4690 1015
rect -4540 1035 -4510 1040
rect -4540 1015 -4535 1035
rect -4535 1015 -4515 1035
rect -4515 1015 -4510 1035
rect -4540 1010 -4510 1015
rect -4360 1035 -4330 1040
rect -4360 1015 -4355 1035
rect -4355 1015 -4335 1035
rect -4335 1015 -4330 1035
rect -4360 1010 -4330 1015
rect -4180 1035 -4150 1040
rect -4180 1015 -4175 1035
rect -4175 1015 -4155 1035
rect -4155 1015 -4150 1035
rect -4180 1010 -4150 1015
rect -4000 1035 -3970 1040
rect -4000 1015 -3995 1035
rect -3995 1015 -3975 1035
rect -3975 1015 -3970 1035
rect -4000 1010 -3970 1015
rect -3820 1035 -3790 1040
rect -3820 1015 -3815 1035
rect -3815 1015 -3795 1035
rect -3795 1015 -3790 1035
rect -3820 1010 -3790 1015
rect -3640 1035 -3610 1040
rect -3640 1015 -3635 1035
rect -3635 1015 -3615 1035
rect -3615 1015 -3610 1035
rect -3640 1010 -3610 1015
rect -3460 1035 -3430 1040
rect -3460 1015 -3455 1035
rect -3455 1015 -3435 1035
rect -3435 1015 -3430 1035
rect -3460 1010 -3430 1015
rect -3280 1035 -3250 1040
rect -3280 1015 -3275 1035
rect -3275 1015 -3255 1035
rect -3255 1015 -3250 1035
rect -3280 1010 -3250 1015
rect -3100 1035 -3070 1040
rect -3100 1015 -3095 1035
rect -3095 1015 -3075 1035
rect -3075 1015 -3070 1035
rect -3100 1010 -3070 1015
rect -2920 1035 -2890 1040
rect -2920 1015 -2915 1035
rect -2915 1015 -2895 1035
rect -2895 1015 -2890 1035
rect -2920 1010 -2890 1015
rect -2740 1035 -2710 1040
rect -2740 1015 -2735 1035
rect -2735 1015 -2715 1035
rect -2715 1015 -2710 1035
rect -2740 1010 -2710 1015
rect -2560 1035 -2530 1040
rect -2560 1015 -2555 1035
rect -2555 1015 -2535 1035
rect -2535 1015 -2530 1035
rect -2560 1010 -2530 1015
rect -2380 1035 -2350 1040
rect -2380 1015 -2375 1035
rect -2375 1015 -2355 1035
rect -2355 1015 -2350 1035
rect -2380 1010 -2350 1015
rect -2200 1035 -2170 1040
rect -2200 1015 -2195 1035
rect -2195 1015 -2175 1035
rect -2175 1015 -2170 1035
rect -2200 1010 -2170 1015
rect -2020 1035 -1990 1040
rect -2020 1015 -2015 1035
rect -2015 1015 -1995 1035
rect -1995 1015 -1990 1035
rect -2020 1010 -1990 1015
rect -1840 1035 -1810 1040
rect -1840 1015 -1835 1035
rect -1835 1015 -1815 1035
rect -1815 1015 -1810 1035
rect -1840 1010 -1810 1015
rect -1660 1035 -1630 1040
rect -1660 1015 -1655 1035
rect -1655 1015 -1635 1035
rect -1635 1015 -1630 1035
rect -1660 1010 -1630 1015
rect -1480 1035 -1450 1040
rect -1480 1015 -1475 1035
rect -1475 1015 -1455 1035
rect -1455 1015 -1450 1035
rect -1480 1010 -1450 1015
rect -1300 1035 -1270 1040
rect -1300 1015 -1295 1035
rect -1295 1015 -1275 1035
rect -1275 1015 -1270 1035
rect -1300 1010 -1270 1015
rect -1120 1035 -1090 1040
rect -1120 1015 -1115 1035
rect -1115 1015 -1095 1035
rect -1095 1015 -1090 1035
rect -1120 1010 -1090 1015
rect -940 1035 -910 1040
rect -940 1015 -935 1035
rect -935 1015 -915 1035
rect -915 1015 -910 1035
rect -940 1010 -910 1015
rect -760 1035 -730 1040
rect -760 1015 -755 1035
rect -755 1015 -735 1035
rect -735 1015 -730 1035
rect -760 1010 -730 1015
rect -10840 980 -10810 985
rect -10840 960 -10835 980
rect -10835 960 -10815 980
rect -10815 960 -10810 980
rect -10840 955 -10810 960
rect -10660 980 -10630 985
rect -10660 960 -10655 980
rect -10655 960 -10635 980
rect -10635 960 -10630 980
rect -10660 955 -10630 960
rect -10480 980 -10450 985
rect -10480 960 -10475 980
rect -10475 960 -10455 980
rect -10455 960 -10450 980
rect -10480 955 -10450 960
rect -10300 980 -10270 985
rect -10300 960 -10295 980
rect -10295 960 -10275 980
rect -10275 960 -10270 980
rect -10300 955 -10270 960
rect -10120 980 -10090 985
rect -10120 960 -10115 980
rect -10115 960 -10095 980
rect -10095 960 -10090 980
rect -10120 955 -10090 960
rect -9940 980 -9910 985
rect -9940 960 -9935 980
rect -9935 960 -9915 980
rect -9915 960 -9910 980
rect -9940 955 -9910 960
rect -9760 980 -9730 985
rect -9760 960 -9755 980
rect -9755 960 -9735 980
rect -9735 960 -9730 980
rect -9760 955 -9730 960
rect -9580 980 -9550 985
rect -9580 960 -9575 980
rect -9575 960 -9555 980
rect -9555 960 -9550 980
rect -9580 955 -9550 960
rect -9400 980 -9370 985
rect -9400 960 -9395 980
rect -9395 960 -9375 980
rect -9375 960 -9370 980
rect -9400 955 -9370 960
rect -9220 980 -9190 985
rect -9220 960 -9215 980
rect -9215 960 -9195 980
rect -9195 960 -9190 980
rect -9220 955 -9190 960
rect -9040 980 -9010 985
rect -9040 960 -9035 980
rect -9035 960 -9015 980
rect -9015 960 -9010 980
rect -9040 955 -9010 960
rect -8860 980 -8830 985
rect -8860 960 -8855 980
rect -8855 960 -8835 980
rect -8835 960 -8830 980
rect -8860 955 -8830 960
rect -8680 980 -8650 985
rect -8680 960 -8675 980
rect -8675 960 -8655 980
rect -8655 960 -8650 980
rect -8680 955 -8650 960
rect -8500 980 -8470 985
rect -8500 960 -8495 980
rect -8495 960 -8475 980
rect -8475 960 -8470 980
rect -8500 955 -8470 960
rect -8320 980 -8290 985
rect -8320 960 -8315 980
rect -8315 960 -8295 980
rect -8295 960 -8290 980
rect -8320 955 -8290 960
rect -8140 980 -8110 985
rect -8140 960 -8135 980
rect -8135 960 -8115 980
rect -8115 960 -8110 980
rect -8140 955 -8110 960
rect -7960 980 -7930 985
rect -7960 960 -7955 980
rect -7955 960 -7935 980
rect -7935 960 -7930 980
rect -7960 955 -7930 960
rect -7780 980 -7750 985
rect -7780 960 -7775 980
rect -7775 960 -7755 980
rect -7755 960 -7750 980
rect -7780 955 -7750 960
rect -7600 980 -7570 985
rect -7600 960 -7595 980
rect -7595 960 -7575 980
rect -7575 960 -7570 980
rect -7600 955 -7570 960
rect -7420 980 -7390 985
rect -7420 960 -7415 980
rect -7415 960 -7395 980
rect -7395 960 -7390 980
rect -7420 955 -7390 960
rect -7240 980 -7210 985
rect -7240 960 -7235 980
rect -7235 960 -7215 980
rect -7215 960 -7210 980
rect -7240 955 -7210 960
rect -7060 980 -7030 985
rect -7060 960 -7055 980
rect -7055 960 -7035 980
rect -7035 960 -7030 980
rect -7060 955 -7030 960
rect -6880 980 -6850 985
rect -6880 960 -6875 980
rect -6875 960 -6855 980
rect -6855 960 -6850 980
rect -6880 955 -6850 960
rect -6700 980 -6670 985
rect -6700 960 -6695 980
rect -6695 960 -6675 980
rect -6675 960 -6670 980
rect -6700 955 -6670 960
rect -6520 980 -6490 985
rect -6520 960 -6515 980
rect -6515 960 -6495 980
rect -6495 960 -6490 980
rect -6520 955 -6490 960
rect -6340 980 -6310 985
rect -6340 960 -6335 980
rect -6335 960 -6315 980
rect -6315 960 -6310 980
rect -6340 955 -6310 960
rect -6160 980 -6130 985
rect -6160 960 -6155 980
rect -6155 960 -6135 980
rect -6135 960 -6130 980
rect -6160 955 -6130 960
rect -5980 980 -5950 985
rect -5980 960 -5975 980
rect -5975 960 -5955 980
rect -5955 960 -5950 980
rect -5980 955 -5950 960
rect -5800 980 -5770 985
rect -5800 960 -5795 980
rect -5795 960 -5775 980
rect -5775 960 -5770 980
rect -5800 955 -5770 960
rect -5620 980 -5590 985
rect -5620 960 -5615 980
rect -5615 960 -5595 980
rect -5595 960 -5590 980
rect -5620 955 -5590 960
rect -5440 980 -5410 985
rect -5440 960 -5435 980
rect -5435 960 -5415 980
rect -5415 960 -5410 980
rect -5440 955 -5410 960
rect -5260 980 -5230 985
rect -5260 960 -5255 980
rect -5255 960 -5235 980
rect -5235 960 -5230 980
rect -5260 955 -5230 960
rect -5080 980 -5050 985
rect -5080 960 -5075 980
rect -5075 960 -5055 980
rect -5055 960 -5050 980
rect -5080 955 -5050 960
rect -4900 980 -4870 985
rect -4900 960 -4895 980
rect -4895 960 -4875 980
rect -4875 960 -4870 980
rect -4900 955 -4870 960
rect -4720 980 -4690 985
rect -4720 960 -4715 980
rect -4715 960 -4695 980
rect -4695 960 -4690 980
rect -4720 955 -4690 960
rect -4540 980 -4510 985
rect -4540 960 -4535 980
rect -4535 960 -4515 980
rect -4515 960 -4510 980
rect -4540 955 -4510 960
rect -4360 980 -4330 985
rect -4360 960 -4355 980
rect -4355 960 -4335 980
rect -4335 960 -4330 980
rect -4360 955 -4330 960
rect -4180 980 -4150 985
rect -4180 960 -4175 980
rect -4175 960 -4155 980
rect -4155 960 -4150 980
rect -4180 955 -4150 960
rect -4000 980 -3970 985
rect -4000 960 -3995 980
rect -3995 960 -3975 980
rect -3975 960 -3970 980
rect -4000 955 -3970 960
rect -3820 980 -3790 985
rect -3820 960 -3815 980
rect -3815 960 -3795 980
rect -3795 960 -3790 980
rect -3820 955 -3790 960
rect -3640 980 -3610 985
rect -3640 960 -3635 980
rect -3635 960 -3615 980
rect -3615 960 -3610 980
rect -3640 955 -3610 960
rect -3460 980 -3430 985
rect -3460 960 -3455 980
rect -3455 960 -3435 980
rect -3435 960 -3430 980
rect -3460 955 -3430 960
rect -3280 980 -3250 985
rect -3280 960 -3275 980
rect -3275 960 -3255 980
rect -3255 960 -3250 980
rect -3280 955 -3250 960
rect -3100 980 -3070 985
rect -3100 960 -3095 980
rect -3095 960 -3075 980
rect -3075 960 -3070 980
rect -3100 955 -3070 960
rect -2920 980 -2890 985
rect -2920 960 -2915 980
rect -2915 960 -2895 980
rect -2895 960 -2890 980
rect -2920 955 -2890 960
rect -2740 980 -2710 985
rect -2740 960 -2735 980
rect -2735 960 -2715 980
rect -2715 960 -2710 980
rect -2740 955 -2710 960
rect -2560 980 -2530 985
rect -2560 960 -2555 980
rect -2555 960 -2535 980
rect -2535 960 -2530 980
rect -2560 955 -2530 960
rect -2380 980 -2350 985
rect -2380 960 -2375 980
rect -2375 960 -2355 980
rect -2355 960 -2350 980
rect -2380 955 -2350 960
rect -2200 980 -2170 985
rect -2200 960 -2195 980
rect -2195 960 -2175 980
rect -2175 960 -2170 980
rect -2200 955 -2170 960
rect -2020 980 -1990 985
rect -2020 960 -2015 980
rect -2015 960 -1995 980
rect -1995 960 -1990 980
rect -2020 955 -1990 960
rect -1840 980 -1810 985
rect -1840 960 -1835 980
rect -1835 960 -1815 980
rect -1815 960 -1810 980
rect -1840 955 -1810 960
rect -1660 980 -1630 985
rect -1660 960 -1655 980
rect -1655 960 -1635 980
rect -1635 960 -1630 980
rect -1660 955 -1630 960
rect -1480 980 -1450 985
rect -1480 960 -1475 980
rect -1475 960 -1455 980
rect -1455 960 -1450 980
rect -1480 955 -1450 960
rect -1300 980 -1270 985
rect -1300 960 -1295 980
rect -1295 960 -1275 980
rect -1275 960 -1270 980
rect -1300 955 -1270 960
rect -1120 980 -1090 985
rect -1120 960 -1115 980
rect -1115 960 -1095 980
rect -1095 960 -1090 980
rect -1120 955 -1090 960
rect -940 980 -910 985
rect -940 960 -935 980
rect -935 960 -915 980
rect -915 960 -910 980
rect -940 955 -910 960
rect -760 980 -730 985
rect -760 960 -755 980
rect -755 960 -735 980
rect -735 960 -730 980
rect -760 955 -730 960
rect -40 1035 -10 1040
rect -40 1015 -35 1035
rect -35 1015 -15 1035
rect -15 1015 -10 1035
rect -40 1010 -10 1015
rect -40 980 -10 985
rect -40 960 -35 980
rect -35 960 -15 980
rect -15 960 -10 980
rect -40 955 -10 960
rect -11695 20 -11665 25
rect -11695 0 -11690 20
rect -11690 0 -11670 20
rect -11670 0 -11665 20
rect -11695 -5 -11665 0
rect -11560 20 -11530 25
rect -11560 0 -11555 20
rect -11555 0 -11535 20
rect -11535 0 -11530 20
rect -11560 -5 -11530 0
rect -10840 20 -10810 25
rect -10840 0 -10835 20
rect -10835 0 -10815 20
rect -10815 0 -10810 20
rect -10840 -5 -10810 0
rect -10660 20 -10630 25
rect -10660 0 -10655 20
rect -10655 0 -10635 20
rect -10635 0 -10630 20
rect -10660 -5 -10630 0
rect -10480 20 -10450 25
rect -10480 0 -10475 20
rect -10475 0 -10455 20
rect -10455 0 -10450 20
rect -10480 -5 -10450 0
rect -10300 20 -10270 25
rect -10300 0 -10295 20
rect -10295 0 -10275 20
rect -10275 0 -10270 20
rect -10300 -5 -10270 0
rect -10120 20 -10090 25
rect -10120 0 -10115 20
rect -10115 0 -10095 20
rect -10095 0 -10090 20
rect -10120 -5 -10090 0
rect -9940 20 -9910 25
rect -9940 0 -9935 20
rect -9935 0 -9915 20
rect -9915 0 -9910 20
rect -9940 -5 -9910 0
rect -9760 20 -9730 25
rect -9760 0 -9755 20
rect -9755 0 -9735 20
rect -9735 0 -9730 20
rect -9760 -5 -9730 0
rect -9580 20 -9550 25
rect -9580 0 -9575 20
rect -9575 0 -9555 20
rect -9555 0 -9550 20
rect -9580 -5 -9550 0
rect -9400 20 -9370 25
rect -9400 0 -9395 20
rect -9395 0 -9375 20
rect -9375 0 -9370 20
rect -9400 -5 -9370 0
rect -9220 20 -9190 25
rect -9220 0 -9215 20
rect -9215 0 -9195 20
rect -9195 0 -9190 20
rect -9220 -5 -9190 0
rect -9040 20 -9010 25
rect -9040 0 -9035 20
rect -9035 0 -9015 20
rect -9015 0 -9010 20
rect -9040 -5 -9010 0
rect -8860 20 -8830 25
rect -8860 0 -8855 20
rect -8855 0 -8835 20
rect -8835 0 -8830 20
rect -8860 -5 -8830 0
rect -8680 20 -8650 25
rect -8680 0 -8675 20
rect -8675 0 -8655 20
rect -8655 0 -8650 20
rect -8680 -5 -8650 0
rect -8500 20 -8470 25
rect -8500 0 -8495 20
rect -8495 0 -8475 20
rect -8475 0 -8470 20
rect -8500 -5 -8470 0
rect -8320 20 -8290 25
rect -8320 0 -8315 20
rect -8315 0 -8295 20
rect -8295 0 -8290 20
rect -8320 -5 -8290 0
rect -8140 20 -8110 25
rect -8140 0 -8135 20
rect -8135 0 -8115 20
rect -8115 0 -8110 20
rect -8140 -5 -8110 0
rect -7960 20 -7930 25
rect -7960 0 -7955 20
rect -7955 0 -7935 20
rect -7935 0 -7930 20
rect -7960 -5 -7930 0
rect -7780 20 -7750 25
rect -7780 0 -7775 20
rect -7775 0 -7755 20
rect -7755 0 -7750 20
rect -7780 -5 -7750 0
rect -7600 20 -7570 25
rect -7600 0 -7595 20
rect -7595 0 -7575 20
rect -7575 0 -7570 20
rect -7600 -5 -7570 0
rect -7420 20 -7390 25
rect -7420 0 -7415 20
rect -7415 0 -7395 20
rect -7395 0 -7390 20
rect -7420 -5 -7390 0
rect -7240 20 -7210 25
rect -7240 0 -7235 20
rect -7235 0 -7215 20
rect -7215 0 -7210 20
rect -7240 -5 -7210 0
rect -7060 20 -7030 25
rect -7060 0 -7055 20
rect -7055 0 -7035 20
rect -7035 0 -7030 20
rect -7060 -5 -7030 0
rect -6880 20 -6850 25
rect -6880 0 -6875 20
rect -6875 0 -6855 20
rect -6855 0 -6850 20
rect -6880 -5 -6850 0
rect -6700 20 -6670 25
rect -6700 0 -6695 20
rect -6695 0 -6675 20
rect -6675 0 -6670 20
rect -6700 -5 -6670 0
rect -6520 20 -6490 25
rect -6520 0 -6515 20
rect -6515 0 -6495 20
rect -6495 0 -6490 20
rect -6520 -5 -6490 0
rect -6340 20 -6310 25
rect -6340 0 -6335 20
rect -6335 0 -6315 20
rect -6315 0 -6310 20
rect -6340 -5 -6310 0
rect -6160 20 -6130 25
rect -6160 0 -6155 20
rect -6155 0 -6135 20
rect -6135 0 -6130 20
rect -6160 -5 -6130 0
rect -5980 20 -5950 25
rect -5980 0 -5975 20
rect -5975 0 -5955 20
rect -5955 0 -5950 20
rect -5980 -5 -5950 0
rect -5800 20 -5770 25
rect -5800 0 -5795 20
rect -5795 0 -5775 20
rect -5775 0 -5770 20
rect -5800 -5 -5770 0
rect -5620 20 -5590 25
rect -5620 0 -5615 20
rect -5615 0 -5595 20
rect -5595 0 -5590 20
rect -5620 -5 -5590 0
rect -5440 20 -5410 25
rect -5440 0 -5435 20
rect -5435 0 -5415 20
rect -5415 0 -5410 20
rect -5440 -5 -5410 0
rect -5260 20 -5230 25
rect -5260 0 -5255 20
rect -5255 0 -5235 20
rect -5235 0 -5230 20
rect -5260 -5 -5230 0
rect -5080 20 -5050 25
rect -5080 0 -5075 20
rect -5075 0 -5055 20
rect -5055 0 -5050 20
rect -5080 -5 -5050 0
rect -4900 20 -4870 25
rect -4900 0 -4895 20
rect -4895 0 -4875 20
rect -4875 0 -4870 20
rect -4900 -5 -4870 0
rect -4720 20 -4690 25
rect -4720 0 -4715 20
rect -4715 0 -4695 20
rect -4695 0 -4690 20
rect -4720 -5 -4690 0
rect -4540 20 -4510 25
rect -4540 0 -4535 20
rect -4535 0 -4515 20
rect -4515 0 -4510 20
rect -4540 -5 -4510 0
rect -4360 20 -4330 25
rect -4360 0 -4355 20
rect -4355 0 -4335 20
rect -4335 0 -4330 20
rect -4360 -5 -4330 0
rect -4180 20 -4150 25
rect -4180 0 -4175 20
rect -4175 0 -4155 20
rect -4155 0 -4150 20
rect -4180 -5 -4150 0
rect -4000 20 -3970 25
rect -4000 0 -3995 20
rect -3995 0 -3975 20
rect -3975 0 -3970 20
rect -4000 -5 -3970 0
rect -3820 20 -3790 25
rect -3820 0 -3815 20
rect -3815 0 -3795 20
rect -3795 0 -3790 20
rect -3820 -5 -3790 0
rect -3640 20 -3610 25
rect -3640 0 -3635 20
rect -3635 0 -3615 20
rect -3615 0 -3610 20
rect -3640 -5 -3610 0
rect -3460 20 -3430 25
rect -3460 0 -3455 20
rect -3455 0 -3435 20
rect -3435 0 -3430 20
rect -3460 -5 -3430 0
rect -3280 20 -3250 25
rect -3280 0 -3275 20
rect -3275 0 -3255 20
rect -3255 0 -3250 20
rect -3280 -5 -3250 0
rect -3100 20 -3070 25
rect -3100 0 -3095 20
rect -3095 0 -3075 20
rect -3075 0 -3070 20
rect -3100 -5 -3070 0
rect -2920 20 -2890 25
rect -2920 0 -2915 20
rect -2915 0 -2895 20
rect -2895 0 -2890 20
rect -2920 -5 -2890 0
rect -2740 20 -2710 25
rect -2740 0 -2735 20
rect -2735 0 -2715 20
rect -2715 0 -2710 20
rect -2740 -5 -2710 0
rect -2560 20 -2530 25
rect -2560 0 -2555 20
rect -2555 0 -2535 20
rect -2535 0 -2530 20
rect -2560 -5 -2530 0
rect -2380 20 -2350 25
rect -2380 0 -2375 20
rect -2375 0 -2355 20
rect -2355 0 -2350 20
rect -2380 -5 -2350 0
rect -2200 20 -2170 25
rect -2200 0 -2195 20
rect -2195 0 -2175 20
rect -2175 0 -2170 20
rect -2200 -5 -2170 0
rect -2020 20 -1990 25
rect -2020 0 -2015 20
rect -2015 0 -1995 20
rect -1995 0 -1990 20
rect -2020 -5 -1990 0
rect -1840 20 -1810 25
rect -1840 0 -1835 20
rect -1835 0 -1815 20
rect -1815 0 -1810 20
rect -1840 -5 -1810 0
rect -1660 20 -1630 25
rect -1660 0 -1655 20
rect -1655 0 -1635 20
rect -1635 0 -1630 20
rect -1660 -5 -1630 0
rect -1480 20 -1450 25
rect -1480 0 -1475 20
rect -1475 0 -1455 20
rect -1455 0 -1450 20
rect -1480 -5 -1450 0
rect -1300 20 -1270 25
rect -1300 0 -1295 20
rect -1295 0 -1275 20
rect -1275 0 -1270 20
rect -1300 -5 -1270 0
rect -1120 20 -1090 25
rect -1120 0 -1115 20
rect -1115 0 -1095 20
rect -1095 0 -1090 20
rect -1120 -5 -1090 0
rect -940 20 -910 25
rect -940 0 -935 20
rect -935 0 -915 20
rect -915 0 -910 20
rect -940 -5 -910 0
rect -760 20 -730 25
rect -760 0 -755 20
rect -755 0 -735 20
rect -735 0 -730 20
rect -760 -5 -730 0
rect -40 20 -10 25
rect -40 0 -35 20
rect -35 0 -15 20
rect -15 0 -10 20
rect -40 -5 -10 0
rect 95 20 125 25
rect 95 0 100 20
rect 100 0 120 20
rect 120 0 125 20
rect 95 -5 125 0
<< metal2 >>
rect -11700 2000 130 2005
rect -11700 1970 -11695 2000
rect -11665 1970 -11560 2000
rect -11530 1970 -10840 2000
rect -10810 1970 -10660 2000
rect -10630 1970 -10480 2000
rect -10450 1970 -10300 2000
rect -10270 1970 -10120 2000
rect -10090 1970 -9940 2000
rect -9910 1970 -9760 2000
rect -9730 1970 -9580 2000
rect -9550 1970 -9400 2000
rect -9370 1970 -9220 2000
rect -9190 1970 -9040 2000
rect -9010 1970 -8860 2000
rect -8830 1970 -8680 2000
rect -8650 1970 -8500 2000
rect -8470 1970 -8320 2000
rect -8290 1970 -8140 2000
rect -8110 1970 -7960 2000
rect -7930 1970 -7780 2000
rect -7750 1970 -7600 2000
rect -7570 1970 -7420 2000
rect -7390 1970 -7240 2000
rect -7210 1970 -7060 2000
rect -7030 1970 -6880 2000
rect -6850 1970 -6700 2000
rect -6670 1970 -6520 2000
rect -6490 1970 -6340 2000
rect -6310 1970 -6160 2000
rect -6130 1970 -5980 2000
rect -5950 1970 -5800 2000
rect -5770 1970 -5620 2000
rect -5590 1970 -5440 2000
rect -5410 1970 -5260 2000
rect -5230 1970 -5080 2000
rect -5050 1970 -4900 2000
rect -4870 1970 -4720 2000
rect -4690 1970 -4540 2000
rect -4510 1970 -4360 2000
rect -4330 1970 -4180 2000
rect -4150 1970 -4000 2000
rect -3970 1970 -3820 2000
rect -3790 1970 -3640 2000
rect -3610 1970 -3460 2000
rect -3430 1970 -3280 2000
rect -3250 1970 -3100 2000
rect -3070 1970 -2920 2000
rect -2890 1970 -2740 2000
rect -2710 1970 -2560 2000
rect -2530 1970 -2380 2000
rect -2350 1970 -2200 2000
rect -2170 1970 -2020 2000
rect -1990 1970 -1840 2000
rect -1810 1970 -1660 2000
rect -1630 1970 -1480 2000
rect -1450 1970 -1300 2000
rect -1270 1970 -1120 2000
rect -1090 1970 -940 2000
rect -910 1970 -760 2000
rect -730 1970 -40 2000
rect -10 1970 95 2000
rect 125 1970 130 2000
rect -11700 1965 130 1970
rect -11570 1040 -5 1045
rect -11570 1010 -11560 1040
rect -11530 1010 -10840 1040
rect -10810 1010 -10660 1040
rect -10630 1010 -10480 1040
rect -10450 1010 -10300 1040
rect -10270 1010 -10120 1040
rect -10090 1010 -9940 1040
rect -9910 1010 -9760 1040
rect -9730 1010 -9580 1040
rect -9550 1010 -9400 1040
rect -9370 1010 -9220 1040
rect -9190 1010 -9040 1040
rect -9010 1010 -8860 1040
rect -8830 1010 -8680 1040
rect -8650 1010 -8500 1040
rect -8470 1010 -8320 1040
rect -8290 1010 -8140 1040
rect -8110 1010 -7960 1040
rect -7930 1010 -7780 1040
rect -7750 1010 -7600 1040
rect -7570 1010 -7420 1040
rect -7390 1010 -7240 1040
rect -7210 1010 -7060 1040
rect -7030 1010 -6880 1040
rect -6850 1010 -6700 1040
rect -6670 1010 -6520 1040
rect -6490 1010 -6340 1040
rect -6310 1010 -6160 1040
rect -6130 1010 -5980 1040
rect -5950 1010 -5800 1040
rect -5770 1010 -5620 1040
rect -5590 1010 -5440 1040
rect -5410 1010 -5260 1040
rect -5230 1010 -5080 1040
rect -5050 1010 -4900 1040
rect -4870 1010 -4720 1040
rect -4690 1010 -4540 1040
rect -4510 1010 -4360 1040
rect -4330 1010 -4180 1040
rect -4150 1010 -4000 1040
rect -3970 1010 -3820 1040
rect -3790 1010 -3640 1040
rect -3610 1010 -3460 1040
rect -3430 1010 -3280 1040
rect -3250 1010 -3100 1040
rect -3070 1010 -2920 1040
rect -2890 1010 -2740 1040
rect -2710 1010 -2560 1040
rect -2530 1010 -2380 1040
rect -2350 1010 -2200 1040
rect -2170 1010 -2020 1040
rect -1990 1010 -1840 1040
rect -1810 1010 -1660 1040
rect -1630 1010 -1480 1040
rect -1450 1010 -1300 1040
rect -1270 1010 -1120 1040
rect -1090 1010 -940 1040
rect -910 1010 -760 1040
rect -730 1010 -40 1040
rect -10 1010 -5 1040
rect -11570 1005 -5 1010
rect -11565 985 0 990
rect -11565 955 -11560 985
rect -11530 955 -10840 985
rect -10810 955 -10660 985
rect -10630 955 -10480 985
rect -10450 955 -10300 985
rect -10270 955 -10120 985
rect -10090 955 -9940 985
rect -9910 955 -9760 985
rect -9730 955 -9580 985
rect -9550 955 -9400 985
rect -9370 955 -9220 985
rect -9190 955 -9040 985
rect -9010 955 -8860 985
rect -8830 955 -8680 985
rect -8650 955 -8500 985
rect -8470 955 -8320 985
rect -8290 955 -8140 985
rect -8110 955 -7960 985
rect -7930 955 -7780 985
rect -7750 955 -7600 985
rect -7570 955 -7420 985
rect -7390 955 -7240 985
rect -7210 955 -7060 985
rect -7030 955 -6880 985
rect -6850 955 -6700 985
rect -6670 955 -6520 985
rect -6490 955 -6340 985
rect -6310 955 -6160 985
rect -6130 955 -5980 985
rect -5950 955 -5800 985
rect -5770 955 -5620 985
rect -5590 955 -5440 985
rect -5410 955 -5260 985
rect -5230 955 -5080 985
rect -5050 955 -4900 985
rect -4870 955 -4720 985
rect -4690 955 -4540 985
rect -4510 955 -4360 985
rect -4330 955 -4180 985
rect -4150 955 -4000 985
rect -3970 955 -3820 985
rect -3790 955 -3640 985
rect -3610 955 -3460 985
rect -3430 955 -3280 985
rect -3250 955 -3100 985
rect -3070 955 -2920 985
rect -2890 955 -2740 985
rect -2710 955 -2560 985
rect -2530 955 -2380 985
rect -2350 955 -2200 985
rect -2170 955 -2020 985
rect -1990 955 -1840 985
rect -1810 955 -1660 985
rect -1630 955 -1480 985
rect -1450 955 -1300 985
rect -1270 955 -1120 985
rect -1090 955 -940 985
rect -910 955 -760 985
rect -730 955 -40 985
rect -10 955 0 985
rect -11565 950 0 955
rect -11700 25 130 30
rect -11700 -5 -11695 25
rect -11665 -5 -11560 25
rect -11530 -5 -10840 25
rect -10810 -5 -10660 25
rect -10630 -5 -10480 25
rect -10450 -5 -10300 25
rect -10270 -5 -10120 25
rect -10090 -5 -9940 25
rect -9910 -5 -9760 25
rect -9730 -5 -9580 25
rect -9550 -5 -9400 25
rect -9370 -5 -9220 25
rect -9190 -5 -9040 25
rect -9010 -5 -8860 25
rect -8830 -5 -8680 25
rect -8650 -5 -8500 25
rect -8470 -5 -8320 25
rect -8290 -5 -8140 25
rect -8110 -5 -7960 25
rect -7930 -5 -7780 25
rect -7750 -5 -7600 25
rect -7570 -5 -7420 25
rect -7390 -5 -7240 25
rect -7210 -5 -7060 25
rect -7030 -5 -6880 25
rect -6850 -5 -6700 25
rect -6670 -5 -6520 25
rect -6490 -5 -6340 25
rect -6310 -5 -6160 25
rect -6130 -5 -5980 25
rect -5950 -5 -5800 25
rect -5770 -5 -5620 25
rect -5590 -5 -5440 25
rect -5410 -5 -5260 25
rect -5230 -5 -5080 25
rect -5050 -5 -4900 25
rect -4870 -5 -4720 25
rect -4690 -5 -4540 25
rect -4510 -5 -4360 25
rect -4330 -5 -4180 25
rect -4150 -5 -4000 25
rect -3970 -5 -3820 25
rect -3790 -5 -3640 25
rect -3610 -5 -3460 25
rect -3430 -5 -3280 25
rect -3250 -5 -3100 25
rect -3070 -5 -2920 25
rect -2890 -5 -2740 25
rect -2710 -5 -2560 25
rect -2530 -5 -2380 25
rect -2350 -5 -2200 25
rect -2170 -5 -2020 25
rect -1990 -5 -1840 25
rect -1810 -5 -1660 25
rect -1630 -5 -1480 25
rect -1450 -5 -1300 25
rect -1270 -5 -1120 25
rect -1090 -5 -940 25
rect -910 -5 -760 25
rect -730 -5 -40 25
rect -10 -5 95 25
rect 125 -5 130 25
rect -11700 -10 130 -5
<< labels >>
rlabel metal2 -11560 970 -11560 970 1 VDDA
port 1 n
rlabel metal2 -11560 10 -11560 10 1 VSSA
port 2 n
rlabel locali -11555 710 -11555 710 1 X
rlabel locali -11555 630 -11555 630 1 P1
port 3 n
rlabel locali -11555 590 -11555 590 1 P2
port 4 n
rlabel locali -11555 310 -11555 310 1 N2
port 5 n
rlabel locali -11555 270 -11555 270 1 N1
port 6 n
rlabel locali -11555 550 -11555 550 1 Z
rlabel locali -11555 430 -11555 430 1 INP
port 7 n
rlabel locali -11555 470 -11555 470 1 INM
port 8 n
rlabel locali -11555 510 -11555 510 1 OUT
port 9 n
rlabel locali -11555 350 -11555 350 1 YP
rlabel locali -11555 390 -11555 390 1 YM
rlabel metal2 -10 1025 -10 1025 5 VDDA
port 1 n
rlabel metal2 -10 1985 -10 1985 5 VSSA
port 2 n
<< end >>
